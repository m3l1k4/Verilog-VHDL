//`timescale 1ns / 1ps
module test_bench_lab_5();


reg clk_tb, rst_tb,CLOCK_50_tb;

wire  [4:0] lfsr_tb;
wire out_sync_tb;
logic [11:0] sino_tb, mod_sig_tb ;
logic out_sync_sig;
logic Clock_1KHz;
logic [11:0] modulated_signal;

wire [4:0] lf_out;

assign modulated_signal = out_sync_sig*sino_tb;

LFSR lfsr_tbr(
.Clock_1KHz(Clock_1KHz),
.rst(rst_tb),
.lfsr_out(lfsr_tb)

);


// for testing remove after
Generate_Arbitrary_Divided_Clk32 
clk_1Hz
(
.inclk(CLOCK_50_tb),
.outclk(Clock_1KHz), //Clock_1KHz
.outclk_Not(),
.div_clk_count(5),  // 1hz 32'h17D7840
.Reset(rst_tb)); 




edge_detect detec_tb( 

// receiveing sub ssytem
.clk_receive(CLOCK_50_tb),
.reset(rst_tb),
.out_edge(out_sync_sig), // synnced signal
// sending subsys
.clk_send(Clock_1KHz), // lfsr clock
.en(lfsr_tb[0])  //lfsr zeroth bit


);




/*
 sig_mod_2 mood_tb(
//input clock,
//input reset,
//.sync_sig(out_sync),
.lfsr_0(out_sync_tb),
.org_wave(sino_tb),
.mod_sig(mod_sig_tb)

);
		
	
		
waveform_gen waves_tb(

 // -- system signals
  .clk(CLOCK_50_tb),       //  : in  std_logic;
  .reset(!rst_tb),     //  : in  std_logic;
  
 // -- clock-enable
 .en(1'b1),         // : in  std_logic;
  
  //-- NCO frequency control
 .phase_inc(258),   //inc = Fout⋅232/ Fs 0.5   //(3e-6(2^32))/50 + 0.5  = 258.19803776 =258   3hz
  
//  -- Output waveforms
  .sin_out(sino_tb),   // 
  .cos_out(),   //  
  .squ_out(),  //   
  .saw_out() );  //  	
*/		
//*/
initial forever begin
// slow clock
clk_tb = 1;
#5;
clk_tb = 0;
#5;

end 

initial forever begin
// fast clock
CLOCK_50_tb = 1;
#1;
CLOCK_50_tb = 0;
#1;
end

initial begin

rst_tb = 1;
#1;
rst_tb = 0;
#1;
rst_tb = 1;
#1;
rst_tb = 0;
#1;

end


initial forever begin

sino_tb=12'h000;#1; sino_tb=12'h003;#1; sino_tb=12'h006;#1; sino_tb=12'h009;#1; sino_tb=12'h00d;#1; sino_tb=12'h010;#1; sino_tb=12'h013;#1; sino_tb=12'h016;#1; 
sino_tb=12'h019;#1; sino_tb=12'h01c;#1; sino_tb=12'h01f;#1; sino_tb=12'h023;#1; sino_tb=12'h026;#1; sino_tb=12'h029;#1; sino_tb=12'h02c;#1; sino_tb=12'h02f;#1; 
sino_tb=12'h032;#1; sino_tb=12'h035;#1; sino_tb=12'h039;#1; sino_tb=12'h03c;#1; sino_tb=12'h03f;#1; sino_tb=12'h042;#1; sino_tb=12'h045;#1; sino_tb=12'h048;#1; 
sino_tb=12'h04b;#1; sino_tb=12'h04e;#1; sino_tb=12'h052;#1; sino_tb=12'h055;#1; sino_tb=12'h058;#1; sino_tb=12'h05b;#1; sino_tb=12'h05e;#1; sino_tb=12'h061;#1; 
sino_tb=12'h064;#1; sino_tb=12'h068;#1; sino_tb=12'h06b;#1; sino_tb=12'h06e;#1; sino_tb=12'h071;#1; sino_tb=12'h074;#1; sino_tb=12'h077;#1; sino_tb=12'h07a;#1; 
sino_tb=12'h07e;#1; sino_tb=12'h081;#1; sino_tb=12'h084;#1; sino_tb=12'h087;#1; sino_tb=12'h08a;#1; sino_tb=12'h08d;#1; sino_tb=12'h090;#1; sino_tb=12'h093;#1; 
sino_tb=12'h097;#1; sino_tb=12'h09a;#1; sino_tb=12'h09d;#1; sino_tb=12'h0a0;#1; sino_tb=12'h0a3;#1; sino_tb=12'h0a6;#1; sino_tb=12'h0a9;#1; sino_tb=12'h0ac;#1; 
sino_tb=12'h0b0;#1; sino_tb=12'h0b3;#1; sino_tb=12'h0b6;#1; sino_tb=12'h0b9;#1; sino_tb=12'h0bc;#1; sino_tb=12'h0bf;#1; sino_tb=12'h0c2;#1; sino_tb=12'h0c6;#1; 
sino_tb=12'h0c9;#1; sino_tb=12'h0cc;#1; sino_tb=12'h0cf;#1; sino_tb=12'h0d2;#1; sino_tb=12'h0d5;#1; sino_tb=12'h0d8;#1; sino_tb=12'h0db;#1; sino_tb=12'h0df;#1; 
sino_tb=12'h0e2;#1; sino_tb=12'h0e5;#1; sino_tb=12'h0e8;#1; sino_tb=12'h0eb;#1; sino_tb=12'h0ee;#1; sino_tb=12'h0f1;#1; sino_tb=12'h0f4;#1; sino_tb=12'h0f7;#1; 
sino_tb=12'h0fb;#1; sino_tb=12'h0fe;#1; sino_tb=12'h101;#1; sino_tb=12'h104;#1; sino_tb=12'h107;#1; sino_tb=12'h10a;#1; sino_tb=12'h10d;#1; sino_tb=12'h110;#1; 
sino_tb=12'h113;#1; sino_tb=12'h117;#1; sino_tb=12'h11a;#1; sino_tb=12'h11d;#1; sino_tb=12'h120;#1; sino_tb=12'h123;#1; sino_tb=12'h126;#1; sino_tb=12'h129;#1; 
sino_tb=12'h12c;#1; sino_tb=12'h12f;#1; sino_tb=12'h133;#1; sino_tb=12'h136;#1; sino_tb=12'h139;#1; sino_tb=12'h13c;#1; sino_tb=12'h13f;#1; sino_tb=12'h142;#1; 
sino_tb=12'h145;#1; sino_tb=12'h148;#1; sino_tb=12'h14b;#1; sino_tb=12'h14e;#1; sino_tb=12'h152;#1; sino_tb=12'h155;#1; sino_tb=12'h158;#1; sino_tb=12'h15b;#1; 
sino_tb=12'h15e;#1; sino_tb=12'h161;#1; sino_tb=12'h164;#1; sino_tb=12'h167;#1; sino_tb=12'h16a;#1; sino_tb=12'h16d;#1; sino_tb=12'h171;#1; sino_tb=12'h174;#1; 
sino_tb=12'h177;#1; sino_tb=12'h17a;#1; sino_tb=12'h17d;#1; sino_tb=12'h180;#1; sino_tb=12'h183;#1; sino_tb=12'h186;#1; sino_tb=12'h189;#1; sino_tb=12'h18c;#1; 
sino_tb=12'h18f;#1; sino_tb=12'h192;#1; sino_tb=12'h196;#1; sino_tb=12'h199;#1; sino_tb=12'h19c;#1; sino_tb=12'h19f;#1; sino_tb=12'h1a2;#1; sino_tb=12'h1a5;#1; 
sino_tb=12'h1a8;#1; sino_tb=12'h1ab;#1; sino_tb=12'h1ae;#1; sino_tb=12'h1b1;#1; sino_tb=12'h1b4;#1; sino_tb=12'h1b7;#1; sino_tb=12'h1ba;#1; sino_tb=12'h1bd;#1; 
sino_tb=12'h1c1;#1; sino_tb=12'h1c4;#1; sino_tb=12'h1c7;#1; sino_tb=12'h1ca;#1; sino_tb=12'h1cd;#1; sino_tb=12'h1d0;#1; sino_tb=12'h1d3;#1; sino_tb=12'h1d6;#1; 
sino_tb=12'h1d9;#1; sino_tb=12'h1dc;#1; sino_tb=12'h1df;#1; sino_tb=12'h1e2;#1; sino_tb=12'h1e5;#1; sino_tb=12'h1e8;#1; sino_tb=12'h1eb;#1; sino_tb=12'h1ee;#1; 
sino_tb=12'h1f1;#1; sino_tb=12'h1f4;#1; sino_tb=12'h1f7;#1; sino_tb=12'h1fb;#1; sino_tb=12'h1fe;#1; sino_tb=12'h201;#1; sino_tb=12'h204;#1; sino_tb=12'h207;#1; 
sino_tb=12'h20a;#1; sino_tb=12'h20d;#1; sino_tb=12'h210;#1; sino_tb=12'h213;#1; sino_tb=12'h216;#1; sino_tb=12'h219;#1; sino_tb=12'h21c;#1; sino_tb=12'h21f;#1; 
sino_tb=12'h222;#1; sino_tb=12'h225;#1; sino_tb=12'h228;#1; sino_tb=12'h22b;#1; sino_tb=12'h22e;#1; sino_tb=12'h231;#1; sino_tb=12'h234;#1; sino_tb=12'h237;#1; 
sino_tb=12'h23a;#1; sino_tb=12'h23d;#1; sino_tb=12'h240;#1; sino_tb=12'h243;#1; sino_tb=12'h246;#1; sino_tb=12'h249;#1; sino_tb=12'h24c;#1; sino_tb=12'h24f;#1; 
sino_tb=12'h252;#1; sino_tb=12'h255;#1; sino_tb=12'h258;#1; sino_tb=12'h25b;#1; sino_tb=12'h25e;#1; sino_tb=12'h261;#1; sino_tb=12'h264;#1; sino_tb=12'h267;#1; 
sino_tb=12'h26a;#1; sino_tb=12'h26d;#1; sino_tb=12'h270;#1; sino_tb=12'h273;#1; sino_tb=12'h276;#1; sino_tb=12'h279;#1; sino_tb=12'h27c;#1; sino_tb=12'h27f;#1; 
sino_tb=12'h282;#1; sino_tb=12'h285;#1; sino_tb=12'h288;#1; sino_tb=12'h28b;#1; sino_tb=12'h28e;#1; sino_tb=12'h291;#1; sino_tb=12'h294;#1; sino_tb=12'h297;#1; 
sino_tb=12'h29a;#1; sino_tb=12'h29d;#1; sino_tb=12'h2a0;#1; sino_tb=12'h2a3;#1; sino_tb=12'h2a6;#1; sino_tb=12'h2a9;#1; sino_tb=12'h2ac;#1; sino_tb=12'h2af;#1; 
sino_tb=12'h2b2;#1; sino_tb=12'h2b5;#1; sino_tb=12'h2b8;#1; sino_tb=12'h2ba;#1; sino_tb=12'h2bd;#1; sino_tb=12'h2c0;#1; sino_tb=12'h2c3;#1; sino_tb=12'h2c6;#1; 
sino_tb=12'h2c9;#1; sino_tb=12'h2cc;#1; sino_tb=12'h2cf;#1; sino_tb=12'h2d2;#1; sino_tb=12'h2d5;#1; sino_tb=12'h2d8;#1; sino_tb=12'h2db;#1; sino_tb=12'h2de;#1; 
sino_tb=12'h2e1;#1; sino_tb=12'h2e4;#1; sino_tb=12'h2e7;#1; sino_tb=12'h2e9;#1; sino_tb=12'h2ec;#1; sino_tb=12'h2ef;#1; sino_tb=12'h2f2;#1; sino_tb=12'h2f5;#1; 
sino_tb=12'h2f8;#1; sino_tb=12'h2fb;#1; sino_tb=12'h2fe;#1; sino_tb=12'h301;#1; sino_tb=12'h304;#1; sino_tb=12'h307;#1; sino_tb=12'h30a;#1; sino_tb=12'h30c;#1; 
sino_tb=12'h30f;#1; sino_tb=12'h312;#1; sino_tb=12'h315;#1; sino_tb=12'h318;#1; sino_tb=12'h31b;#1; sino_tb=12'h31e;#1; sino_tb=12'h321;#1; sino_tb=12'h324;#1; 
sino_tb=12'h327;#1; sino_tb=12'h329;#1; sino_tb=12'h32c;#1; sino_tb=12'h32f;#1; sino_tb=12'h332;#1; sino_tb=12'h335;#1; sino_tb=12'h338;#1; sino_tb=12'h33b;#1; 
sino_tb=12'h33e;#1; sino_tb=12'h340;#1; sino_tb=12'h343;#1; sino_tb=12'h346;#1; sino_tb=12'h349;#1; sino_tb=12'h34c;#1; sino_tb=12'h34f;#1; sino_tb=12'h352;#1; 
sino_tb=12'h354;#1; sino_tb=12'h357;#1; sino_tb=12'h35a;#1; sino_tb=12'h35d;#1; sino_tb=12'h360;#1; sino_tb=12'h363;#1; sino_tb=12'h366;#1; sino_tb=12'h368;#1; 
sino_tb=12'h36b;#1; sino_tb=12'h36e;#1; sino_tb=12'h371;#1; sino_tb=12'h374;#1; sino_tb=12'h377;#1; sino_tb=12'h379;#1; sino_tb=12'h37c;#1; sino_tb=12'h37f;#1; 
sino_tb=12'h382;#1; sino_tb=12'h385;#1; sino_tb=12'h387;#1; sino_tb=12'h38a;#1; sino_tb=12'h38d;#1; sino_tb=12'h390;#1; sino_tb=12'h393;#1; sino_tb=12'h396;#1; 
sino_tb=12'h398;#1; sino_tb=12'h39b;#1; sino_tb=12'h39e;#1; sino_tb=12'h3a1;#1; sino_tb=12'h3a4;#1; sino_tb=12'h3a6;#1; sino_tb=12'h3a9;#1; sino_tb=12'h3ac;#1; 
sino_tb=12'h3af;#1; sino_tb=12'h3b2;#1; sino_tb=12'h3b4;#1; sino_tb=12'h3b7;#1; sino_tb=12'h3ba;#1; sino_tb=12'h3bd;#1; sino_tb=12'h3bf;#1; sino_tb=12'h3c2;#1; 
sino_tb=12'h3c5;#1; sino_tb=12'h3c8;#1; sino_tb=12'h3ca;#1; sino_tb=12'h3cd;#1; sino_tb=12'h3d0;#1; sino_tb=12'h3d3;#1; sino_tb=12'h3d6;#1; sino_tb=12'h3d8;#1; 
sino_tb=12'h3db;#1; sino_tb=12'h3de;#1; sino_tb=12'h3e1;#1; sino_tb=12'h3e3;#1; sino_tb=12'h3e6;#1; sino_tb=12'h3e9;#1; sino_tb=12'h3eb;#1; sino_tb=12'h3ee;#1; 
sino_tb=12'h3f1;#1; sino_tb=12'h3f4;#1; sino_tb=12'h3f6;#1; sino_tb=12'h3f9;#1; sino_tb=12'h3fc;#1; sino_tb=12'h3ff;#1; sino_tb=12'h401;#1; sino_tb=12'h404;#1; 
sino_tb=12'h407;#1; sino_tb=12'h409;#1; sino_tb=12'h40c;#1; sino_tb=12'h40f;#1; sino_tb=12'h412;#1; sino_tb=12'h414;#1; sino_tb=12'h417;#1; sino_tb=12'h41a;#1; 
sino_tb=12'h41c;#1; sino_tb=12'h41f;#1; sino_tb=12'h422;#1; sino_tb=12'h424;#1; sino_tb=12'h427;#1; sino_tb=12'h42a;#1; sino_tb=12'h42c;#1; sino_tb=12'h42f;#1; 
sino_tb=12'h432;#1; sino_tb=12'h435;#1; sino_tb=12'h437;#1; sino_tb=12'h43a;#1; sino_tb=12'h43d;#1; sino_tb=12'h43f;#1; sino_tb=12'h442;#1; sino_tb=12'h444;#1; 
sino_tb=12'h447;#1; sino_tb=12'h44a;#1; sino_tb=12'h44c;#1; sino_tb=12'h44f;#1; sino_tb=12'h452;#1; sino_tb=12'h454;#1; sino_tb=12'h457;#1; sino_tb=12'h45a;#1; 
sino_tb=12'h45c;#1; sino_tb=12'h45f;#1; sino_tb=12'h462;#1; sino_tb=12'h464;#1; sino_tb=12'h467;#1; sino_tb=12'h469;#1; sino_tb=12'h46c;#1; sino_tb=12'h46f;#1; 
sino_tb=12'h471;#1; sino_tb=12'h474;#1; sino_tb=12'h476;#1; sino_tb=12'h479;#1; sino_tb=12'h47c;#1; sino_tb=12'h47e;#1; sino_tb=12'h481;#1; sino_tb=12'h483;#1; 
sino_tb=12'h486;#1; sino_tb=12'h489;#1; sino_tb=12'h48b;#1; sino_tb=12'h48e;#1; sino_tb=12'h490;#1; sino_tb=12'h493;#1; sino_tb=12'h496;#1; sino_tb=12'h498;#1; 
sino_tb=12'h49b;#1; sino_tb=12'h49d;#1; sino_tb=12'h4a0;#1; sino_tb=12'h4a2;#1; sino_tb=12'h4a5;#1; sino_tb=12'h4a7;#1; sino_tb=12'h4aa;#1; sino_tb=12'h4ad;#1; 
sino_tb=12'h4af;#1; sino_tb=12'h4b2;#1; sino_tb=12'h4b4;#1; sino_tb=12'h4b7;#1; sino_tb=12'h4b9;#1; sino_tb=12'h4bc;#1; sino_tb=12'h4be;#1; sino_tb=12'h4c1;#1; 
sino_tb=12'h4c3;#1; sino_tb=12'h4c6;#1; sino_tb=12'h4c8;#1; sino_tb=12'h4cb;#1; sino_tb=12'h4cd;#1; sino_tb=12'h4d0;#1; sino_tb=12'h4d2;#1; sino_tb=12'h4d5;#1; 
sino_tb=12'h4d7;#1; sino_tb=12'h4da;#1; sino_tb=12'h4dc;#1; sino_tb=12'h4df;#1; sino_tb=12'h4e1;#1; sino_tb=12'h4e4;#1; sino_tb=12'h4e6;#1; sino_tb=12'h4e9;#1; 
sino_tb=12'h4eb;#1; sino_tb=12'h4ee;#1; sino_tb=12'h4f0;#1; sino_tb=12'h4f3;#1; sino_tb=12'h4f5;#1; sino_tb=12'h4f8;#1; sino_tb=12'h4fa;#1; sino_tb=12'h4fd;#1; 
sino_tb=12'h4ff;#1; sino_tb=12'h502;#1; sino_tb=12'h504;#1; sino_tb=12'h506;#1; sino_tb=12'h509;#1; sino_tb=12'h50b;#1; sino_tb=12'h50e;#1; sino_tb=12'h510;#1; 
sino_tb=12'h513;#1; sino_tb=12'h515;#1; sino_tb=12'h517;#1; sino_tb=12'h51a;#1; sino_tb=12'h51c;#1; sino_tb=12'h51f;#1; sino_tb=12'h521;#1; sino_tb=12'h524;#1; 
sino_tb=12'h526;#1; sino_tb=12'h528;#1; sino_tb=12'h52b;#1; sino_tb=12'h52d;#1; sino_tb=12'h530;#1; sino_tb=12'h532;#1; sino_tb=12'h534;#1; sino_tb=12'h537;#1; 
sino_tb=12'h539;#1; sino_tb=12'h53b;#1; sino_tb=12'h53e;#1; sino_tb=12'h540;#1; sino_tb=12'h543;#1; sino_tb=12'h545;#1; sino_tb=12'h547;#1; sino_tb=12'h54a;#1; 
sino_tb=12'h54c;#1; sino_tb=12'h54e;#1; sino_tb=12'h551;#1; sino_tb=12'h553;#1; sino_tb=12'h555;#1; sino_tb=12'h558;#1; sino_tb=12'h55a;#1; sino_tb=12'h55c;#1; 
sino_tb=12'h55f;#1; sino_tb=12'h561;#1; sino_tb=12'h563;#1; sino_tb=12'h566;#1; sino_tb=12'h568;#1; sino_tb=12'h56a;#1; sino_tb=12'h56d;#1; sino_tb=12'h56f;#1; 
sino_tb=12'h571;#1; sino_tb=12'h573;#1; sino_tb=12'h576;#1; sino_tb=12'h578;#1; sino_tb=12'h57a;#1; sino_tb=12'h57d;#1; sino_tb=12'h57f;#1; sino_tb=12'h581;#1; 
sino_tb=12'h583;#1; sino_tb=12'h586;#1; sino_tb=12'h588;#1; sino_tb=12'h58a;#1; sino_tb=12'h58d;#1; sino_tb=12'h58f;#1; sino_tb=12'h591;#1; sino_tb=12'h593;#1; 
sino_tb=12'h596;#1; sino_tb=12'h598;#1; sino_tb=12'h59a;#1; sino_tb=12'h59c;#1; sino_tb=12'h59f;#1; sino_tb=12'h5a1;#1; sino_tb=12'h5a3;#1; sino_tb=12'h5a5;#1; 
sino_tb=12'h5a7;#1; sino_tb=12'h5aa;#1; sino_tb=12'h5ac;#1; sino_tb=12'h5ae;#1; sino_tb=12'h5b0;#1; sino_tb=12'h5b3;#1; sino_tb=12'h5b5;#1; sino_tb=12'h5b7;#1; 
sino_tb=12'h5b9;#1; sino_tb=12'h5bb;#1; sino_tb=12'h5bd;#1; sino_tb=12'h5c0;#1; sino_tb=12'h5c2;#1; sino_tb=12'h5c4;#1; sino_tb=12'h5c6;#1; sino_tb=12'h5c8;#1; 
sino_tb=12'h5cb;#1; sino_tb=12'h5cd;#1; sino_tb=12'h5cf;#1; sino_tb=12'h5d1;#1; sino_tb=12'h5d3;#1; sino_tb=12'h5d5;#1; sino_tb=12'h5d7;#1; sino_tb=12'h5da;#1; 
sino_tb=12'h5dc;#1; sino_tb=12'h5de;#1; sino_tb=12'h5e0;#1; sino_tb=12'h5e2;#1; sino_tb=12'h5e4;#1; sino_tb=12'h5e6;#1; sino_tb=12'h5e9;#1; sino_tb=12'h5eb;#1; 
sino_tb=12'h5ed;#1; sino_tb=12'h5ef;#1; sino_tb=12'h5f1;#1; sino_tb=12'h5f3;#1; sino_tb=12'h5f5;#1; sino_tb=12'h5f7;#1; sino_tb=12'h5f9;#1; sino_tb=12'h5fb;#1; 
sino_tb=12'h5fd;#1; sino_tb=12'h600;#1; sino_tb=12'h602;#1; sino_tb=12'h604;#1; sino_tb=12'h606;#1; sino_tb=12'h608;#1; sino_tb=12'h60a;#1; sino_tb=12'h60c;#1; 
sino_tb=12'h60e;#1; sino_tb=12'h610;#1; sino_tb=12'h612;#1; sino_tb=12'h614;#1; sino_tb=12'h616;#1; sino_tb=12'h618;#1; sino_tb=12'h61a;#1; sino_tb=12'h61c;#1; 
sino_tb=12'h61e;#1; sino_tb=12'h620;#1; sino_tb=12'h622;#1; sino_tb=12'h624;#1; sino_tb=12'h626;#1; sino_tb=12'h628;#1; sino_tb=12'h62a;#1; sino_tb=12'h62c;#1; 
sino_tb=12'h62e;#1; sino_tb=12'h630;#1; sino_tb=12'h632;#1; sino_tb=12'h634;#1; sino_tb=12'h636;#1; sino_tb=12'h638;#1; sino_tb=12'h63a;#1; sino_tb=12'h63c;#1; 
sino_tb=12'h63e;#1; sino_tb=12'h640;#1; sino_tb=12'h642;#1; sino_tb=12'h644;#1; sino_tb=12'h646;#1; sino_tb=12'h648;#1; sino_tb=12'h64a;#1; sino_tb=12'h64c;#1; 
sino_tb=12'h64e;#1; sino_tb=12'h650;#1; sino_tb=12'h652;#1; sino_tb=12'h654;#1; sino_tb=12'h655;#1; sino_tb=12'h657;#1; sino_tb=12'h659;#1; sino_tb=12'h65b;#1; 
sino_tb=12'h65d;#1; sino_tb=12'h65f;#1; sino_tb=12'h661;#1; sino_tb=12'h663;#1; sino_tb=12'h665;#1; sino_tb=12'h667;#1; sino_tb=12'h668;#1; sino_tb=12'h66a;#1; 
sino_tb=12'h66c;#1; sino_tb=12'h66e;#1; sino_tb=12'h670;#1; sino_tb=12'h672;#1; sino_tb=12'h674;#1; sino_tb=12'h675;#1; sino_tb=12'h677;#1; sino_tb=12'h679;#1; 
sino_tb=12'h67b;#1; sino_tb=12'h67d;#1; sino_tb=12'h67f;#1; sino_tb=12'h681;#1; sino_tb=12'h682;#1; sino_tb=12'h684;#1; sino_tb=12'h686;#1; sino_tb=12'h688;#1; 
sino_tb=12'h68a;#1; sino_tb=12'h68b;#1; sino_tb=12'h68d;#1; sino_tb=12'h68f;#1; sino_tb=12'h691;#1; sino_tb=12'h693;#1; sino_tb=12'h694;#1; sino_tb=12'h696;#1; 
sino_tb=12'h698;#1; sino_tb=12'h69a;#1; sino_tb=12'h69b;#1; sino_tb=12'h69d;#1; sino_tb=12'h69f;#1; sino_tb=12'h6a1;#1; sino_tb=12'h6a3;#1; sino_tb=12'h6a4;#1; 
sino_tb=12'h6a6;#1; sino_tb=12'h6a8;#1; sino_tb=12'h6a9;#1; sino_tb=12'h6ab;#1; sino_tb=12'h6ad;#1; sino_tb=12'h6af;#1; sino_tb=12'h6b0;#1; sino_tb=12'h6b2;#1; 
sino_tb=12'h6b4;#1; sino_tb=12'h6b6;#1; sino_tb=12'h6b7;#1; sino_tb=12'h6b9;#1; sino_tb=12'h6bb;#1; sino_tb=12'h6bc;#1; sino_tb=12'h6be;#1; sino_tb=12'h6c0;#1; 
sino_tb=12'h6c1;#1; sino_tb=12'h6c3;#1; sino_tb=12'h6c5;#1; sino_tb=12'h6c6;#1; sino_tb=12'h6c8;#1; sino_tb=12'h6ca;#1; sino_tb=12'h6cb;#1; sino_tb=12'h6cd;#1; 
sino_tb=12'h6cf;#1; sino_tb=12'h6d0;#1; sino_tb=12'h6d2;#1; sino_tb=12'h6d4;#1; sino_tb=12'h6d5;#1; sino_tb=12'h6d7;#1; sino_tb=12'h6d9;#1; sino_tb=12'h6da;#1; 
sino_tb=12'h6dc;#1; sino_tb=12'h6dd;#1; sino_tb=12'h6df;#1; sino_tb=12'h6e1;#1; sino_tb=12'h6e2;#1; sino_tb=12'h6e4;#1; sino_tb=12'h6e5;#1; sino_tb=12'h6e7;#1; 
sino_tb=12'h6e9;#1; sino_tb=12'h6ea;#1; sino_tb=12'h6ec;#1; sino_tb=12'h6ed;#1; sino_tb=12'h6ef;#1; sino_tb=12'h6f0;#1; sino_tb=12'h6f2;#1; sino_tb=12'h6f4;#1; 
sino_tb=12'h6f5;#1; sino_tb=12'h6f7;#1; sino_tb=12'h6f8;#1; sino_tb=12'h6fa;#1; sino_tb=12'h6fb;#1; sino_tb=12'h6fd;#1; sino_tb=12'h6fe;#1; sino_tb=12'h700;#1; 
sino_tb=12'h701;#1; sino_tb=12'h703;#1; sino_tb=12'h704;#1; sino_tb=12'h706;#1; sino_tb=12'h707;#1; sino_tb=12'h709;#1; sino_tb=12'h70a;#1; sino_tb=12'h70c;#1; 
sino_tb=12'h70d;#1; sino_tb=12'h70f;#1; sino_tb=12'h710;#1; sino_tb=12'h712;#1; sino_tb=12'h713;#1; sino_tb=12'h715;#1; sino_tb=12'h716;#1; sino_tb=12'h718;#1; 
sino_tb=12'h719;#1; sino_tb=12'h71a;#1; sino_tb=12'h71c;#1; sino_tb=12'h71d;#1; sino_tb=12'h71f;#1; sino_tb=12'h720;#1; sino_tb=12'h722;#1; sino_tb=12'h723;#1; 
sino_tb=12'h724;#1; sino_tb=12'h726;#1; sino_tb=12'h727;#1; sino_tb=12'h729;#1; sino_tb=12'h72a;#1; sino_tb=12'h72b;#1; sino_tb=12'h72d;#1; sino_tb=12'h72e;#1; 
sino_tb=12'h730;#1; sino_tb=12'h731;#1; sino_tb=12'h732;#1; sino_tb=12'h734;#1; sino_tb=12'h735;#1; sino_tb=12'h736;#1; sino_tb=12'h738;#1; sino_tb=12'h739;#1; 
sino_tb=12'h73a;#1; sino_tb=12'h73c;#1; sino_tb=12'h73d;#1; sino_tb=12'h73e;#1; sino_tb=12'h740;#1; sino_tb=12'h741;#1; sino_tb=12'h742;#1; sino_tb=12'h744;#1; 
sino_tb=12'h745;#1; sino_tb=12'h746;#1; sino_tb=12'h748;#1; sino_tb=12'h749;#1; sino_tb=12'h74a;#1; sino_tb=12'h74c;#1; sino_tb=12'h74d;#1; sino_tb=12'h74e;#1; 
sino_tb=12'h74f;#1; sino_tb=12'h751;#1; sino_tb=12'h752;#1; sino_tb=12'h753;#1; sino_tb=12'h754;#1; sino_tb=12'h756;#1; sino_tb=12'h757;#1; sino_tb=12'h758;#1; 
sino_tb=12'h759;#1; sino_tb=12'h75b;#1; sino_tb=12'h75c;#1; sino_tb=12'h75d;#1; sino_tb=12'h75e;#1; sino_tb=12'h760;#1; sino_tb=12'h761;#1; sino_tb=12'h762;#1; 
sino_tb=12'h763;#1; sino_tb=12'h764;#1; sino_tb=12'h766;#1; sino_tb=12'h767;#1; sino_tb=12'h768;#1; sino_tb=12'h769;#1; sino_tb=12'h76a;#1; sino_tb=12'h76b;#1; 
sino_tb=12'h76d;#1; sino_tb=12'h76e;#1; sino_tb=12'h76f;#1; sino_tb=12'h770;#1; sino_tb=12'h771;#1; sino_tb=12'h772;#1; sino_tb=12'h774;#1; sino_tb=12'h775;#1; 
sino_tb=12'h776;#1; sino_tb=12'h777;#1; sino_tb=12'h778;#1; sino_tb=12'h779;#1; sino_tb=12'h77a;#1; sino_tb=12'h77b;#1; sino_tb=12'h77d;#1; sino_tb=12'h77e;#1; 
sino_tb=12'h77f;#1; sino_tb=12'h780;#1; sino_tb=12'h781;#1; sino_tb=12'h782;#1; sino_tb=12'h783;#1; sino_tb=12'h784;#1; sino_tb=12'h785;#1; sino_tb=12'h786;#1; 
sino_tb=12'h787;#1; sino_tb=12'h788;#1; sino_tb=12'h789;#1; sino_tb=12'h78a;#1; sino_tb=12'h78c;#1; sino_tb=12'h78d;#1; sino_tb=12'h78e;#1; sino_tb=12'h78f;#1; 
sino_tb=12'h790;#1; sino_tb=12'h791;#1; sino_tb=12'h792;#1; sino_tb=12'h793;#1; sino_tb=12'h794;#1; sino_tb=12'h795;#1; sino_tb=12'h796;#1; sino_tb=12'h797;#1; 
sino_tb=12'h798;#1; sino_tb=12'h799;#1; sino_tb=12'h79a;#1; sino_tb=12'h79b;#1; sino_tb=12'h79c;#1; sino_tb=12'h79d;#1; sino_tb=12'h79e;#1; sino_tb=12'h79e;#1; 
sino_tb=12'h79f;#1; sino_tb=12'h7a0;#1; sino_tb=12'h7a1;#1; sino_tb=12'h7a2;#1; sino_tb=12'h7a3;#1; sino_tb=12'h7a4;#1; sino_tb=12'h7a5;#1; sino_tb=12'h7a6;#1; 
sino_tb=12'h7a7;#1; sino_tb=12'h7a8;#1; sino_tb=12'h7a9;#1; sino_tb=12'h7aa;#1; sino_tb=12'h7aa;#1; sino_tb=12'h7ab;#1; sino_tb=12'h7ac;#1; sino_tb=12'h7ad;#1; 
sino_tb=12'h7ae;#1; sino_tb=12'h7af;#1; sino_tb=12'h7b0;#1; sino_tb=12'h7b1;#1; sino_tb=12'h7b1;#1; sino_tb=12'h7b2;#1; sino_tb=12'h7b3;#1; sino_tb=12'h7b4;#1; 
sino_tb=12'h7b5;#1; sino_tb=12'h7b6;#1; sino_tb=12'h7b7;#1; sino_tb=12'h7b7;#1; sino_tb=12'h7b8;#1; sino_tb=12'h7b9;#1; sino_tb=12'h7ba;#1; sino_tb=12'h7bb;#1; 
sino_tb=12'h7bb;#1; sino_tb=12'h7bc;#1; sino_tb=12'h7bd;#1; sino_tb=12'h7be;#1; sino_tb=12'h7bf;#1; sino_tb=12'h7bf;#1; sino_tb=12'h7c0;#1; sino_tb=12'h7c1;#1; 
sino_tb=12'h7c2;#1; sino_tb=12'h7c2;#1; sino_tb=12'h7c3;#1; sino_tb=12'h7c4;#1; sino_tb=12'h7c5;#1; sino_tb=12'h7c5;#1; sino_tb=12'h7c6;#1; sino_tb=12'h7c7;#1; 
sino_tb=12'h7c8;#1; sino_tb=12'h7c8;#1; sino_tb=12'h7c9;#1; sino_tb=12'h7ca;#1; sino_tb=12'h7ca;#1; sino_tb=12'h7cb;#1; sino_tb=12'h7cc;#1; sino_tb=12'h7cd;#1; 
sino_tb=12'h7cd;#1; sino_tb=12'h7ce;#1; sino_tb=12'h7cf;#1; sino_tb=12'h7cf;#1; sino_tb=12'h7d0;#1; sino_tb=12'h7d1;#1; sino_tb=12'h7d1;#1; sino_tb=12'h7d2;#1; 
sino_tb=12'h7d3;#1; sino_tb=12'h7d3;#1; sino_tb=12'h7d4;#1; sino_tb=12'h7d5;#1; sino_tb=12'h7d5;#1; sino_tb=12'h7d6;#1; sino_tb=12'h7d6;#1; sino_tb=12'h7d7;#1; 
sino_tb=12'h7d8;#1; sino_tb=12'h7d8;#1; sino_tb=12'h7d9;#1; sino_tb=12'h7d9;#1; sino_tb=12'h7da;#1; sino_tb=12'h7db;#1; sino_tb=12'h7db;#1; sino_tb=12'h7dc;#1; 
sino_tb=12'h7dc;#1; sino_tb=12'h7dd;#1; sino_tb=12'h7de;#1; sino_tb=12'h7de;#1; sino_tb=12'h7df;#1; sino_tb=12'h7df;#1; sino_tb=12'h7e0;#1; sino_tb=12'h7e0;#1; 
sino_tb=12'h7e1;#1; sino_tb=12'h7e1;#1; sino_tb=12'h7e2;#1; sino_tb=12'h7e2;#1; sino_tb=12'h7e3;#1; sino_tb=12'h7e3;#1; sino_tb=12'h7e4;#1; sino_tb=12'h7e5;#1; 
sino_tb=12'h7e5;#1; sino_tb=12'h7e6;#1; sino_tb=12'h7e6;#1; sino_tb=12'h7e6;#1; sino_tb=12'h7e7;#1; sino_tb=12'h7e7;#1; sino_tb=12'h7e8;#1; sino_tb=12'h7e8;#1; 
sino_tb=12'h7e9;#1; sino_tb=12'h7e9;#1; sino_tb=12'h7ea;#1; sino_tb=12'h7ea;#1; sino_tb=12'h7eb;#1; sino_tb=12'h7eb;#1; sino_tb=12'h7ec;#1; sino_tb=12'h7ec;#1; 
sino_tb=12'h7ec;#1; sino_tb=12'h7ed;#1; sino_tb=12'h7ed;#1; sino_tb=12'h7ee;#1; sino_tb=12'h7ee;#1; sino_tb=12'h7ee;#1; sino_tb=12'h7ef;#1; sino_tb=12'h7ef;#1; 
sino_tb=12'h7f0;#1; sino_tb=12'h7f0;#1; sino_tb=12'h7f0;#1; sino_tb=12'h7f1;#1; sino_tb=12'h7f1;#1; sino_tb=12'h7f1;#1; sino_tb=12'h7f2;#1; sino_tb=12'h7f2;#1; 
sino_tb=12'h7f3;#1; sino_tb=12'h7f3;#1; sino_tb=12'h7f3;#1; sino_tb=12'h7f4;#1; sino_tb=12'h7f4;#1; sino_tb=12'h7f4;#1; sino_tb=12'h7f5;#1; sino_tb=12'h7f5;#1; 
sino_tb=12'h7f5;#1; sino_tb=12'h7f5;#1; sino_tb=12'h7f6;#1; sino_tb=12'h7f6;#1; sino_tb=12'h7f6;#1; sino_tb=12'h7f7;#1; sino_tb=12'h7f7;#1; sino_tb=12'h7f7;#1; 
sino_tb=12'h7f7;#1; sino_tb=12'h7f8;#1; sino_tb=12'h7f8;#1; sino_tb=12'h7f8;#1; sino_tb=12'h7f8;#1; sino_tb=12'h7f9;#1; sino_tb=12'h7f9;#1; sino_tb=12'h7f9;#1; 
sino_tb=12'h7f9;#1; sino_tb=12'h7fa;#1; sino_tb=12'h7fa;#1; sino_tb=12'h7fa;#1; sino_tb=12'h7fa;#1; sino_tb=12'h7fb;#1; sino_tb=12'h7fb;#1; sino_tb=12'h7fb;#1; 
sino_tb=12'h7fb;#1; sino_tb=12'h7fb;#1; sino_tb=12'h7fc;#1; sino_tb=12'h7fc;#1; sino_tb=12'h7fc;#1; sino_tb=12'h7fc;#1; sino_tb=12'h7fc;#1; sino_tb=12'h7fc;#1; 
sino_tb=12'h7fd;#1; sino_tb=12'h7fd;#1; sino_tb=12'h7fd;#1; sino_tb=12'h7fd;#1; sino_tb=12'h7fd;#1; sino_tb=12'h7fd;#1; sino_tb=12'h7fd;#1; sino_tb=12'h7fd;#1; 
sino_tb=12'h7fe;#1; sino_tb=12'h7fe;#1; sino_tb=12'h7fe;#1; sino_tb=12'h7fe;#1; sino_tb=12'h7fe;#1; sino_tb=12'h7fe;#1; sino_tb=12'h7fe;#1; sino_tb=12'h7fe;#1; 
sino_tb=12'h7fe;#1; sino_tb=12'h7fe;#1; sino_tb=12'h7ff;#1; sino_tb=12'h7ff;#1; sino_tb=12'h7ff;#1; sino_tb=12'h7ff;#1; sino_tb=12'h7ff;#1; sino_tb=12'h7ff;#1; 
sino_tb=12'h7ff;#1; sino_tb=12'h7ff;#1; sino_tb=12'h7ff;#1; sino_tb=12'h7ff;#1; sino_tb=12'h7ff;#1; sino_tb=12'h7ff;#1; sino_tb=12'h7ff;#1; sino_tb=12'h7ff;#1; 
sino_tb=12'h7ff;#1; sino_tb=12'h7ff;#1; sino_tb=12'h7ff;#1; sino_tb=12'h7ff;#1; sino_tb=12'h7ff;#1; sino_tb=12'h7ff;#1; sino_tb=12'h7ff;#1; sino_tb=12'h7ff;#1; 
sino_tb=12'h7ff;#1; sino_tb=12'h7ff;#1; sino_tb=12'h7ff;#1; sino_tb=12'h7ff;#1; sino_tb=12'h7ff;#1; sino_tb=12'h7ff;#1; sino_tb=12'h7ff;#1; sino_tb=12'h7fe;#1; 
sino_tb=12'h7fe;#1; sino_tb=12'h7fe;#1; sino_tb=12'h7fe;#1; sino_tb=12'h7fe;#1; sino_tb=12'h7fe;#1; sino_tb=12'h7fe;#1; sino_tb=12'h7fe;#1; sino_tb=12'h7fe;#1; 
sino_tb=12'h7fe;#1; sino_tb=12'h7fd;#1; sino_tb=12'h7fd;#1; sino_tb=12'h7fd;#1; sino_tb=12'h7fd;#1; sino_tb=12'h7fd;#1; sino_tb=12'h7fd;#1; sino_tb=12'h7fd;#1; 
sino_tb=12'h7fd;#1; sino_tb=12'h7fc;#1; sino_tb=12'h7fc;#1; sino_tb=12'h7fc;#1; sino_tb=12'h7fc;#1; sino_tb=12'h7fc;#1; sino_tb=12'h7fc;#1; sino_tb=12'h7fb;#1; 
sino_tb=12'h7fb;#1; sino_tb=12'h7fb;#1; sino_tb=12'h7fb;#1; sino_tb=12'h7fb;#1; sino_tb=12'h7fa;#1; sino_tb=12'h7fa;#1; sino_tb=12'h7fa;#1; sino_tb=12'h7fa;#1; 
sino_tb=12'h7f9;#1; sino_tb=12'h7f9;#1; sino_tb=12'h7f9;#1; sino_tb=12'h7f9;#1; sino_tb=12'h7f8;#1; sino_tb=12'h7f8;#1; sino_tb=12'h7f8;#1; sino_tb=12'h7f8;#1; 
sino_tb=12'h7f7;#1; sino_tb=12'h7f7;#1; sino_tb=12'h7f7;#1; sino_tb=12'h7f7;#1; sino_tb=12'h7f6;#1; sino_tb=12'h7f6;#1; sino_tb=12'h7f6;#1; sino_tb=12'h7f5;#1; 
sino_tb=12'h7f5;#1; sino_tb=12'h7f5;#1; sino_tb=12'h7f5;#1; sino_tb=12'h7f4;#1; sino_tb=12'h7f4;#1; sino_tb=12'h7f4;#1; sino_tb=12'h7f3;#1; sino_tb=12'h7f3;#1; 
sino_tb=12'h7f3;#1; sino_tb=12'h7f2;#1; sino_tb=12'h7f2;#1; sino_tb=12'h7f1;#1; sino_tb=12'h7f1;#1; sino_tb=12'h7f1;#1; sino_tb=12'h7f0;#1; sino_tb=12'h7f0;#1; 
sino_tb=12'h7f0;#1; sino_tb=12'h7ef;#1; sino_tb=12'h7ef;#1; sino_tb=12'h7ee;#1; sino_tb=12'h7ee;#1; sino_tb=12'h7ee;#1; sino_tb=12'h7ed;#1; sino_tb=12'h7ed;#1; 
sino_tb=12'h7ec;#1; sino_tb=12'h7ec;#1; sino_tb=12'h7ec;#1; sino_tb=12'h7eb;#1; sino_tb=12'h7eb;#1; sino_tb=12'h7ea;#1; sino_tb=12'h7ea;#1; sino_tb=12'h7e9;#1; 
sino_tb=12'h7e9;#1; sino_tb=12'h7e8;#1; sino_tb=12'h7e8;#1; sino_tb=12'h7e7;#1; sino_tb=12'h7e7;#1; sino_tb=12'h7e6;#1; sino_tb=12'h7e6;#1; sino_tb=12'h7e6;#1; 
sino_tb=12'h7e5;#1; sino_tb=12'h7e5;#1; sino_tb=12'h7e4;#1; sino_tb=12'h7e3;#1; sino_tb=12'h7e3;#1; sino_tb=12'h7e2;#1; sino_tb=12'h7e2;#1; sino_tb=12'h7e1;#1; 
sino_tb=12'h7e1;#1; sino_tb=12'h7e0;#1; sino_tb=12'h7e0;#1; sino_tb=12'h7df;#1; sino_tb=12'h7df;#1; sino_tb=12'h7de;#1; sino_tb=12'h7de;#1; sino_tb=12'h7dd;#1; 
sino_tb=12'h7dc;#1; sino_tb=12'h7dc;#1; sino_tb=12'h7db;#1; sino_tb=12'h7db;#1; sino_tb=12'h7da;#1; sino_tb=12'h7d9;#1; sino_tb=12'h7d9;#1; sino_tb=12'h7d8;#1; 
sino_tb=12'h7d8;#1; sino_tb=12'h7d7;#1; sino_tb=12'h7d6;#1; sino_tb=12'h7d6;#1; sino_tb=12'h7d5;#1; sino_tb=12'h7d5;#1; sino_tb=12'h7d4;#1; sino_tb=12'h7d3;#1; 
sino_tb=12'h7d3;#1; sino_tb=12'h7d2;#1; sino_tb=12'h7d1;#1; sino_tb=12'h7d1;#1; sino_tb=12'h7d0;#1; sino_tb=12'h7cf;#1; sino_tb=12'h7cf;#1; sino_tb=12'h7ce;#1; 
sino_tb=12'h7cd;#1; sino_tb=12'h7cd;#1; sino_tb=12'h7cc;#1; sino_tb=12'h7cb;#1; sino_tb=12'h7ca;#1; sino_tb=12'h7ca;#1; sino_tb=12'h7c9;#1; sino_tb=12'h7c8;#1; 
sino_tb=12'h7c8;#1; sino_tb=12'h7c7;#1; sino_tb=12'h7c6;#1; sino_tb=12'h7c5;#1; sino_tb=12'h7c5;#1; sino_tb=12'h7c4;#1; sino_tb=12'h7c3;#1; sino_tb=12'h7c2;#1; 
sino_tb=12'h7c2;#1; sino_tb=12'h7c1;#1; sino_tb=12'h7c0;#1; sino_tb=12'h7bf;#1; sino_tb=12'h7bf;#1; sino_tb=12'h7be;#1; sino_tb=12'h7bd;#1; sino_tb=12'h7bc;#1; 
sino_tb=12'h7bb;#1; sino_tb=12'h7bb;#1; sino_tb=12'h7ba;#1; sino_tb=12'h7b9;#1; sino_tb=12'h7b8;#1; sino_tb=12'h7b7;#1; sino_tb=12'h7b7;#1; sino_tb=12'h7b6;#1; 
sino_tb=12'h7b5;#1; sino_tb=12'h7b4;#1; sino_tb=12'h7b3;#1; sino_tb=12'h7b2;#1; sino_tb=12'h7b1;#1; sino_tb=12'h7b1;#1; sino_tb=12'h7b0;#1; sino_tb=12'h7af;#1; 
sino_tb=12'h7ae;#1; sino_tb=12'h7ad;#1; sino_tb=12'h7ac;#1; sino_tb=12'h7ab;#1; sino_tb=12'h7aa;#1; sino_tb=12'h7aa;#1; sino_tb=12'h7a9;#1; sino_tb=12'h7a8;#1; 
sino_tb=12'h7a7;#1; sino_tb=12'h7a6;#1; sino_tb=12'h7a5;#1; sino_tb=12'h7a4;#1; sino_tb=12'h7a3;#1; sino_tb=12'h7a2;#1; sino_tb=12'h7a1;#1; sino_tb=12'h7a0;#1; 
sino_tb=12'h79f;#1; sino_tb=12'h79e;#1; sino_tb=12'h79e;#1; sino_tb=12'h79d;#1; sino_tb=12'h79c;#1; sino_tb=12'h79b;#1; sino_tb=12'h79a;#1; sino_tb=12'h799;#1; 
sino_tb=12'h798;#1; sino_tb=12'h797;#1; sino_tb=12'h796;#1; sino_tb=12'h795;#1; sino_tb=12'h794;#1; sino_tb=12'h793;#1; sino_tb=12'h792;#1; sino_tb=12'h791;#1; 
sino_tb=12'h790;#1; sino_tb=12'h78f;#1; sino_tb=12'h78e;#1; sino_tb=12'h78d;#1; sino_tb=12'h78c;#1; sino_tb=12'h78a;#1; sino_tb=12'h789;#1; sino_tb=12'h788;#1; 
sino_tb=12'h787;#1; sino_tb=12'h786;#1; sino_tb=12'h785;#1; sino_tb=12'h784;#1; sino_tb=12'h783;#1; sino_tb=12'h782;#1; sino_tb=12'h781;#1; sino_tb=12'h780;#1; 
sino_tb=12'h77f;#1; sino_tb=12'h77e;#1; sino_tb=12'h77d;#1; sino_tb=12'h77b;#1; sino_tb=12'h77a;#1; sino_tb=12'h779;#1; sino_tb=12'h778;#1; sino_tb=12'h777;#1; 
sino_tb=12'h776;#1; sino_tb=12'h775;#1; sino_tb=12'h774;#1; sino_tb=12'h772;#1; sino_tb=12'h771;#1; sino_tb=12'h770;#1; sino_tb=12'h76f;#1; sino_tb=12'h76e;#1; 
sino_tb=12'h76d;#1; sino_tb=12'h76b;#1; sino_tb=12'h76a;#1; sino_tb=12'h769;#1; sino_tb=12'h768;#1; sino_tb=12'h767;#1; sino_tb=12'h766;#1; sino_tb=12'h764;#1; 
sino_tb=12'h763;#1; sino_tb=12'h762;#1; sino_tb=12'h761;#1; sino_tb=12'h760;#1; sino_tb=12'h75e;#1; sino_tb=12'h75d;#1; sino_tb=12'h75c;#1; sino_tb=12'h75b;#1; 
sino_tb=12'h759;#1; sino_tb=12'h758;#1; sino_tb=12'h757;#1; sino_tb=12'h756;#1; sino_tb=12'h754;#1; sino_tb=12'h753;#1; sino_tb=12'h752;#1; sino_tb=12'h751;#1; 
sino_tb=12'h74f;#1; sino_tb=12'h74e;#1; sino_tb=12'h74d;#1; sino_tb=12'h74c;#1; sino_tb=12'h74a;#1; sino_tb=12'h749;#1; sino_tb=12'h748;#1; sino_tb=12'h746;#1; 
sino_tb=12'h745;#1; sino_tb=12'h744;#1; sino_tb=12'h742;#1; sino_tb=12'h741;#1; sino_tb=12'h740;#1; sino_tb=12'h73e;#1; sino_tb=12'h73d;#1; sino_tb=12'h73c;#1; 
sino_tb=12'h73a;#1; sino_tb=12'h739;#1; sino_tb=12'h738;#1; sino_tb=12'h736;#1; sino_tb=12'h735;#1; sino_tb=12'h734;#1; sino_tb=12'h732;#1; sino_tb=12'h731;#1; 
sino_tb=12'h730;#1; sino_tb=12'h72e;#1; sino_tb=12'h72d;#1; sino_tb=12'h72b;#1; sino_tb=12'h72a;#1; sino_tb=12'h729;#1; sino_tb=12'h727;#1; sino_tb=12'h726;#1; 
sino_tb=12'h724;#1; sino_tb=12'h723;#1; sino_tb=12'h722;#1; sino_tb=12'h720;#1; sino_tb=12'h71f;#1; sino_tb=12'h71d;#1; sino_tb=12'h71c;#1; sino_tb=12'h71a;#1; 
sino_tb=12'h719;#1; sino_tb=12'h718;#1; sino_tb=12'h716;#1; sino_tb=12'h715;#1; sino_tb=12'h713;#1; sino_tb=12'h712;#1; sino_tb=12'h710;#1; sino_tb=12'h70f;#1; 
sino_tb=12'h70d;#1; sino_tb=12'h70c;#1; sino_tb=12'h70a;#1; sino_tb=12'h709;#1; sino_tb=12'h707;#1; sino_tb=12'h706;#1; sino_tb=12'h704;#1; sino_tb=12'h703;#1; 
sino_tb=12'h701;#1; sino_tb=12'h700;#1; sino_tb=12'h6fe;#1; sino_tb=12'h6fd;#1; sino_tb=12'h6fb;#1; sino_tb=12'h6fa;#1; sino_tb=12'h6f8;#1; sino_tb=12'h6f7;#1; 
sino_tb=12'h6f5;#1; sino_tb=12'h6f4;#1; sino_tb=12'h6f2;#1; sino_tb=12'h6f0;#1; sino_tb=12'h6ef;#1; sino_tb=12'h6ed;#1; sino_tb=12'h6ec;#1; sino_tb=12'h6ea;#1; 
sino_tb=12'h6e9;#1; sino_tb=12'h6e7;#1; sino_tb=12'h6e5;#1; sino_tb=12'h6e4;#1; sino_tb=12'h6e2;#1; sino_tb=12'h6e1;#1; sino_tb=12'h6df;#1; sino_tb=12'h6dd;#1; 
sino_tb=12'h6dc;#1; sino_tb=12'h6da;#1; sino_tb=12'h6d9;#1; sino_tb=12'h6d7;#1; sino_tb=12'h6d5;#1; sino_tb=12'h6d4;#1; sino_tb=12'h6d2;#1; sino_tb=12'h6d0;#1; 
sino_tb=12'h6cf;#1; sino_tb=12'h6cd;#1; sino_tb=12'h6cb;#1; sino_tb=12'h6ca;#1; sino_tb=12'h6c8;#1; sino_tb=12'h6c6;#1; sino_tb=12'h6c5;#1; sino_tb=12'h6c3;#1; 
sino_tb=12'h6c1;#1; sino_tb=12'h6c0;#1; sino_tb=12'h6be;#1; sino_tb=12'h6bc;#1; sino_tb=12'h6bb;#1; sino_tb=12'h6b9;#1; sino_tb=12'h6b7;#1; sino_tb=12'h6b6;#1; 
sino_tb=12'h6b4;#1; sino_tb=12'h6b2;#1; sino_tb=12'h6b0;#1; sino_tb=12'h6af;#1; sino_tb=12'h6ad;#1; sino_tb=12'h6ab;#1; sino_tb=12'h6a9;#1; sino_tb=12'h6a8;#1; 
sino_tb=12'h6a6;#1; sino_tb=12'h6a4;#1; sino_tb=12'h6a3;#1; sino_tb=12'h6a1;#1; sino_tb=12'h69f;#1; sino_tb=12'h69d;#1; sino_tb=12'h69b;#1; sino_tb=12'h69a;#1; 
sino_tb=12'h698;#1; sino_tb=12'h696;#1; sino_tb=12'h694;#1; sino_tb=12'h693;#1; sino_tb=12'h691;#1; sino_tb=12'h68f;#1; sino_tb=12'h68d;#1; sino_tb=12'h68b;#1; 
sino_tb=12'h68a;#1; sino_tb=12'h688;#1; sino_tb=12'h686;#1; sino_tb=12'h684;#1; sino_tb=12'h682;#1; sino_tb=12'h681;#1; sino_tb=12'h67f;#1; sino_tb=12'h67d;#1; 
sino_tb=12'h67b;#1; sino_tb=12'h679;#1; sino_tb=12'h677;#1; sino_tb=12'h675;#1; sino_tb=12'h674;#1; sino_tb=12'h672;#1; sino_tb=12'h670;#1; sino_tb=12'h66e;#1; 
sino_tb=12'h66c;#1; sino_tb=12'h66a;#1; sino_tb=12'h668;#1; sino_tb=12'h667;#1; sino_tb=12'h665;#1; sino_tb=12'h663;#1; sino_tb=12'h661;#1; sino_tb=12'h65f;#1; 
sino_tb=12'h65d;#1; sino_tb=12'h65b;#1; sino_tb=12'h659;#1; sino_tb=12'h657;#1; sino_tb=12'h655;#1; sino_tb=12'h654;#1; sino_tb=12'h652;#1; sino_tb=12'h650;#1; 
sino_tb=12'h64e;#1; sino_tb=12'h64c;#1; sino_tb=12'h64a;#1; sino_tb=12'h648;#1; sino_tb=12'h646;#1; sino_tb=12'h644;#1; sino_tb=12'h642;#1; sino_tb=12'h640;#1; 
sino_tb=12'h63e;#1; sino_tb=12'h63c;#1; sino_tb=12'h63a;#1; sino_tb=12'h638;#1; sino_tb=12'h636;#1; sino_tb=12'h634;#1; sino_tb=12'h632;#1; sino_tb=12'h630;#1; 
sino_tb=12'h62e;#1; sino_tb=12'h62c;#1; sino_tb=12'h62a;#1; sino_tb=12'h628;#1; sino_tb=12'h626;#1; sino_tb=12'h624;#1; sino_tb=12'h622;#1; sino_tb=12'h620;#1; 
sino_tb=12'h61e;#1; sino_tb=12'h61c;#1; sino_tb=12'h61a;#1; sino_tb=12'h618;#1; sino_tb=12'h616;#1; sino_tb=12'h614;#1; sino_tb=12'h612;#1; sino_tb=12'h610;#1; 
sino_tb=12'h60e;#1; sino_tb=12'h60c;#1; sino_tb=12'h60a;#1; sino_tb=12'h608;#1; sino_tb=12'h606;#1; sino_tb=12'h604;#1; sino_tb=12'h602;#1; sino_tb=12'h600;#1; 
sino_tb=12'h5fd;#1; sino_tb=12'h5fb;#1; sino_tb=12'h5f9;#1; sino_tb=12'h5f7;#1; sino_tb=12'h5f5;#1; sino_tb=12'h5f3;#1; sino_tb=12'h5f1;#1; sino_tb=12'h5ef;#1; 
sino_tb=12'h5ed;#1; sino_tb=12'h5eb;#1; sino_tb=12'h5e9;#1; sino_tb=12'h5e6;#1; sino_tb=12'h5e4;#1; sino_tb=12'h5e2;#1; sino_tb=12'h5e0;#1; sino_tb=12'h5de;#1; 
sino_tb=12'h5dc;#1; sino_tb=12'h5da;#1; sino_tb=12'h5d7;#1; sino_tb=12'h5d5;#1; sino_tb=12'h5d3;#1; sino_tb=12'h5d1;#1; sino_tb=12'h5cf;#1; sino_tb=12'h5cd;#1; 
sino_tb=12'h5cb;#1; sino_tb=12'h5c8;#1; sino_tb=12'h5c6;#1; sino_tb=12'h5c4;#1; sino_tb=12'h5c2;#1; sino_tb=12'h5c0;#1; sino_tb=12'h5bd;#1; sino_tb=12'h5bb;#1; 
sino_tb=12'h5b9;#1; sino_tb=12'h5b7;#1; sino_tb=12'h5b5;#1; sino_tb=12'h5b3;#1; sino_tb=12'h5b0;#1; sino_tb=12'h5ae;#1; sino_tb=12'h5ac;#1; sino_tb=12'h5aa;#1; 
sino_tb=12'h5a7;#1; sino_tb=12'h5a5;#1; sino_tb=12'h5a3;#1; sino_tb=12'h5a1;#1; sino_tb=12'h59f;#1; sino_tb=12'h59c;#1; sino_tb=12'h59a;#1; sino_tb=12'h598;#1; 
sino_tb=12'h596;#1; sino_tb=12'h593;#1; sino_tb=12'h591;#1; sino_tb=12'h58f;#1; sino_tb=12'h58d;#1; sino_tb=12'h58a;#1; sino_tb=12'h588;#1; sino_tb=12'h586;#1; 
sino_tb=12'h583;#1; sino_tb=12'h581;#1; sino_tb=12'h57f;#1; sino_tb=12'h57d;#1; sino_tb=12'h57a;#1; sino_tb=12'h578;#1; sino_tb=12'h576;#1; sino_tb=12'h573;#1; 
sino_tb=12'h571;#1; sino_tb=12'h56f;#1; sino_tb=12'h56d;#1; sino_tb=12'h56a;#1; sino_tb=12'h568;#1; sino_tb=12'h566;#1; sino_tb=12'h563;#1; sino_tb=12'h561;#1; 
sino_tb=12'h55f;#1; sino_tb=12'h55c;#1; sino_tb=12'h55a;#1; sino_tb=12'h558;#1; sino_tb=12'h555;#1; sino_tb=12'h553;#1; sino_tb=12'h551;#1; sino_tb=12'h54e;#1; 
sino_tb=12'h54c;#1; sino_tb=12'h54a;#1; sino_tb=12'h547;#1; sino_tb=12'h545;#1; sino_tb=12'h543;#1; sino_tb=12'h540;#1; sino_tb=12'h53e;#1; sino_tb=12'h53b;#1; 
sino_tb=12'h539;#1; sino_tb=12'h537;#1; sino_tb=12'h534;#1; sino_tb=12'h532;#1; sino_tb=12'h530;#1; sino_tb=12'h52d;#1; sino_tb=12'h52b;#1; sino_tb=12'h528;#1; 
sino_tb=12'h526;#1; sino_tb=12'h524;#1; sino_tb=12'h521;#1; sino_tb=12'h51f;#1; sino_tb=12'h51c;#1; sino_tb=12'h51a;#1; sino_tb=12'h517;#1; sino_tb=12'h515;#1; 
sino_tb=12'h513;#1; sino_tb=12'h510;#1; sino_tb=12'h50e;#1; sino_tb=12'h50b;#1; sino_tb=12'h509;#1; sino_tb=12'h506;#1; sino_tb=12'h504;#1; sino_tb=12'h502;#1; 
sino_tb=12'h4ff;#1; sino_tb=12'h4fd;#1; sino_tb=12'h4fa;#1; sino_tb=12'h4f8;#1; sino_tb=12'h4f5;#1; sino_tb=12'h4f3;#1; sino_tb=12'h4f0;#1; sino_tb=12'h4ee;#1; 
sino_tb=12'h4eb;#1; sino_tb=12'h4e9;#1; sino_tb=12'h4e6;#1; sino_tb=12'h4e4;#1; sino_tb=12'h4e1;#1; sino_tb=12'h4df;#1; sino_tb=12'h4dc;#1; sino_tb=12'h4da;#1; 
sino_tb=12'h4d7;#1; sino_tb=12'h4d5;#1; sino_tb=12'h4d2;#1; sino_tb=12'h4d0;#1; sino_tb=12'h4cd;#1; sino_tb=12'h4cb;#1; sino_tb=12'h4c8;#1; sino_tb=12'h4c6;#1; 
sino_tb=12'h4c3;#1; sino_tb=12'h4c1;#1; sino_tb=12'h4be;#1; sino_tb=12'h4bc;#1; sino_tb=12'h4b9;#1; sino_tb=12'h4b7;#1; sino_tb=12'h4b4;#1; sino_tb=12'h4b2;#1; 
sino_tb=12'h4af;#1; sino_tb=12'h4ad;#1; sino_tb=12'h4aa;#1; sino_tb=12'h4a7;#1; sino_tb=12'h4a5;#1; sino_tb=12'h4a2;#1; sino_tb=12'h4a0;#1; sino_tb=12'h49d;#1; 
sino_tb=12'h49b;#1; sino_tb=12'h498;#1; sino_tb=12'h496;#1; sino_tb=12'h493;#1; sino_tb=12'h490;#1; sino_tb=12'h48e;#1; sino_tb=12'h48b;#1; sino_tb=12'h489;#1; 
sino_tb=12'h486;#1; sino_tb=12'h483;#1; sino_tb=12'h481;#1; sino_tb=12'h47e;#1; sino_tb=12'h47c;#1; sino_tb=12'h479;#1; sino_tb=12'h476;#1; sino_tb=12'h474;#1; 
sino_tb=12'h471;#1; sino_tb=12'h46f;#1; sino_tb=12'h46c;#1; sino_tb=12'h469;#1; sino_tb=12'h467;#1; sino_tb=12'h464;#1; sino_tb=12'h462;#1; sino_tb=12'h45f;#1; 
sino_tb=12'h45c;#1; sino_tb=12'h45a;#1; sino_tb=12'h457;#1; sino_tb=12'h454;#1; sino_tb=12'h452;#1; sino_tb=12'h44f;#1; sino_tb=12'h44c;#1; sino_tb=12'h44a;#1; 
sino_tb=12'h447;#1; sino_tb=12'h444;#1; sino_tb=12'h442;#1; sino_tb=12'h43f;#1; sino_tb=12'h43d;#1; sino_tb=12'h43a;#1; sino_tb=12'h437;#1; sino_tb=12'h435;#1; 
sino_tb=12'h432;#1; sino_tb=12'h42f;#1; sino_tb=12'h42c;#1; sino_tb=12'h42a;#1; sino_tb=12'h427;#1; sino_tb=12'h424;#1; sino_tb=12'h422;#1; sino_tb=12'h41f;#1; 
sino_tb=12'h41c;#1; sino_tb=12'h41a;#1; sino_tb=12'h417;#1; sino_tb=12'h414;#1; sino_tb=12'h412;#1; sino_tb=12'h40f;#1; sino_tb=12'h40c;#1; sino_tb=12'h409;#1; 
sino_tb=12'h407;#1; sino_tb=12'h404;#1; sino_tb=12'h401;#1; sino_tb=12'h3ff;#1; sino_tb=12'h3fc;#1; sino_tb=12'h3f9;#1; sino_tb=12'h3f6;#1; sino_tb=12'h3f4;#1; 
sino_tb=12'h3f1;#1; sino_tb=12'h3ee;#1; sino_tb=12'h3eb;#1; sino_tb=12'h3e9;#1; sino_tb=12'h3e6;#1; sino_tb=12'h3e3;#1; sino_tb=12'h3e1;#1; sino_tb=12'h3de;#1; 
sino_tb=12'h3db;#1; sino_tb=12'h3d8;#1; sino_tb=12'h3d6;#1; sino_tb=12'h3d3;#1; sino_tb=12'h3d0;#1; sino_tb=12'h3cd;#1; sino_tb=12'h3ca;#1; sino_tb=12'h3c8;#1; 
sino_tb=12'h3c5;#1; sino_tb=12'h3c2;#1; sino_tb=12'h3bf;#1; sino_tb=12'h3bd;#1; sino_tb=12'h3ba;#1; sino_tb=12'h3b7;#1; sino_tb=12'h3b4;#1; sino_tb=12'h3b2;#1; 
sino_tb=12'h3af;#1; sino_tb=12'h3ac;#1; sino_tb=12'h3a9;#1; sino_tb=12'h3a6;#1; sino_tb=12'h3a4;#1; sino_tb=12'h3a1;#1; sino_tb=12'h39e;#1; sino_tb=12'h39b;#1; 
sino_tb=12'h398;#1; sino_tb=12'h396;#1; sino_tb=12'h393;#1; sino_tb=12'h390;#1; sino_tb=12'h38d;#1; sino_tb=12'h38a;#1; sino_tb=12'h387;#1; sino_tb=12'h385;#1; 
sino_tb=12'h382;#1; sino_tb=12'h37f;#1; sino_tb=12'h37c;#1; sino_tb=12'h379;#1; sino_tb=12'h377;#1; sino_tb=12'h374;#1; sino_tb=12'h371;#1; sino_tb=12'h36e;#1; 
sino_tb=12'h36b;#1; sino_tb=12'h368;#1; sino_tb=12'h366;#1; sino_tb=12'h363;#1; sino_tb=12'h360;#1; sino_tb=12'h35d;#1; sino_tb=12'h35a;#1; sino_tb=12'h357;#1; 
sino_tb=12'h354;#1; sino_tb=12'h352;#1; sino_tb=12'h34f;#1; sino_tb=12'h34c;#1; sino_tb=12'h349;#1; sino_tb=12'h346;#1; sino_tb=12'h343;#1; sino_tb=12'h340;#1; 
sino_tb=12'h33e;#1; sino_tb=12'h33b;#1; sino_tb=12'h338;#1; sino_tb=12'h335;#1; sino_tb=12'h332;#1; sino_tb=12'h32f;#1; sino_tb=12'h32c;#1; sino_tb=12'h329;#1; 
sino_tb=12'h327;#1; sino_tb=12'h324;#1; sino_tb=12'h321;#1; sino_tb=12'h31e;#1; sino_tb=12'h31b;#1; sino_tb=12'h318;#1; sino_tb=12'h315;#1; sino_tb=12'h312;#1; 
sino_tb=12'h30f;#1; sino_tb=12'h30c;#1; sino_tb=12'h30a;#1; sino_tb=12'h307;#1; sino_tb=12'h304;#1; sino_tb=12'h301;#1; sino_tb=12'h2fe;#1; sino_tb=12'h2fb;#1; 
sino_tb=12'h2f8;#1; sino_tb=12'h2f5;#1; sino_tb=12'h2f2;#1; sino_tb=12'h2ef;#1; sino_tb=12'h2ec;#1; sino_tb=12'h2e9;#1; sino_tb=12'h2e7;#1; sino_tb=12'h2e4;#1; 
sino_tb=12'h2e1;#1; sino_tb=12'h2de;#1; sino_tb=12'h2db;#1; sino_tb=12'h2d8;#1; sino_tb=12'h2d5;#1; sino_tb=12'h2d2;#1; sino_tb=12'h2cf;#1; sino_tb=12'h2cc;#1; 
sino_tb=12'h2c9;#1; sino_tb=12'h2c6;#1; sino_tb=12'h2c3;#1; sino_tb=12'h2c0;#1; sino_tb=12'h2bd;#1; sino_tb=12'h2ba;#1; sino_tb=12'h2b8;#1; sino_tb=12'h2b5;#1; 
sino_tb=12'h2b2;#1; sino_tb=12'h2af;#1; sino_tb=12'h2ac;#1; sino_tb=12'h2a9;#1; sino_tb=12'h2a6;#1; sino_tb=12'h2a3;#1; sino_tb=12'h2a0;#1; sino_tb=12'h29d;#1; 
sino_tb=12'h29a;#1; sino_tb=12'h297;#1; sino_tb=12'h294;#1; sino_tb=12'h291;#1; sino_tb=12'h28e;#1; sino_tb=12'h28b;#1; sino_tb=12'h288;#1; sino_tb=12'h285;#1; 
sino_tb=12'h282;#1; sino_tb=12'h27f;#1; sino_tb=12'h27c;#1; sino_tb=12'h279;#1; sino_tb=12'h276;#1; sino_tb=12'h273;#1; sino_tb=12'h270;#1; sino_tb=12'h26d;#1; 
sino_tb=12'h26a;#1; sino_tb=12'h267;#1; sino_tb=12'h264;#1; sino_tb=12'h261;#1; sino_tb=12'h25e;#1; sino_tb=12'h25b;#1; sino_tb=12'h258;#1; sino_tb=12'h255;#1; 
sino_tb=12'h252;#1; sino_tb=12'h24f;#1; sino_tb=12'h24c;#1; sino_tb=12'h249;#1; sino_tb=12'h246;#1; sino_tb=12'h243;#1; sino_tb=12'h240;#1; sino_tb=12'h23d;#1; 
sino_tb=12'h23a;#1; sino_tb=12'h237;#1; sino_tb=12'h234;#1; sino_tb=12'h231;#1; sino_tb=12'h22e;#1; sino_tb=12'h22b;#1; sino_tb=12'h228;#1; sino_tb=12'h225;#1; 
sino_tb=12'h222;#1; sino_tb=12'h21f;#1; sino_tb=12'h21c;#1; sino_tb=12'h219;#1; sino_tb=12'h216;#1; sino_tb=12'h213;#1; sino_tb=12'h210;#1; sino_tb=12'h20d;#1; 
sino_tb=12'h20a;#1; sino_tb=12'h207;#1; sino_tb=12'h204;#1; sino_tb=12'h201;#1; sino_tb=12'h1fe;#1; sino_tb=12'h1fb;#1; sino_tb=12'h1f7;#1; sino_tb=12'h1f4;#1; 
sino_tb=12'h1f1;#1; sino_tb=12'h1ee;#1; sino_tb=12'h1eb;#1; sino_tb=12'h1e8;#1; sino_tb=12'h1e5;#1; sino_tb=12'h1e2;#1; sino_tb=12'h1df;#1; sino_tb=12'h1dc;#1; 
sino_tb=12'h1d9;#1; sino_tb=12'h1d6;#1; sino_tb=12'h1d3;#1; sino_tb=12'h1d0;#1; sino_tb=12'h1cd;#1; sino_tb=12'h1ca;#1; sino_tb=12'h1c7;#1; sino_tb=12'h1c4;#1; 
sino_tb=12'h1c1;#1; sino_tb=12'h1bd;#1; sino_tb=12'h1ba;#1; sino_tb=12'h1b7;#1; sino_tb=12'h1b4;#1; sino_tb=12'h1b1;#1; sino_tb=12'h1ae;#1; sino_tb=12'h1ab;#1; 
sino_tb=12'h1a8;#1; sino_tb=12'h1a5;#1; sino_tb=12'h1a2;#1; sino_tb=12'h19f;#1; sino_tb=12'h19c;#1; sino_tb=12'h199;#1; sino_tb=12'h196;#1; sino_tb=12'h192;#1; 
sino_tb=12'h18f;#1; sino_tb=12'h18c;#1; sino_tb=12'h189;#1; sino_tb=12'h186;#1; sino_tb=12'h183;#1; sino_tb=12'h180;#1; sino_tb=12'h17d;#1; sino_tb=12'h17a;#1; 
sino_tb=12'h177;#1; sino_tb=12'h174;#1; sino_tb=12'h171;#1; sino_tb=12'h16d;#1; sino_tb=12'h16a;#1; sino_tb=12'h167;#1; sino_tb=12'h164;#1; sino_tb=12'h161;#1; 
sino_tb=12'h15e;#1; sino_tb=12'h15b;#1; sino_tb=12'h158;#1; sino_tb=12'h155;#1; sino_tb=12'h152;#1; sino_tb=12'h14e;#1; sino_tb=12'h14b;#1; sino_tb=12'h148;#1; 
sino_tb=12'h145;#1; sino_tb=12'h142;#1; sino_tb=12'h13f;#1; sino_tb=12'h13c;#1; sino_tb=12'h139;#1; sino_tb=12'h136;#1; sino_tb=12'h133;#1; sino_tb=12'h12f;#1; 
sino_tb=12'h12c;#1; sino_tb=12'h129;#1; sino_tb=12'h126;#1; sino_tb=12'h123;#1; sino_tb=12'h120;#1; sino_tb=12'h11d;#1; sino_tb=12'h11a;#1; sino_tb=12'h117;#1; 
sino_tb=12'h113;#1; sino_tb=12'h110;#1; sino_tb=12'h10d;#1; sino_tb=12'h10a;#1; sino_tb=12'h107;#1; sino_tb=12'h104;#1; sino_tb=12'h101;#1; sino_tb=12'h0fe;#1; 
sino_tb=12'h0fb;#1; sino_tb=12'h0f7;#1; sino_tb=12'h0f4;#1; sino_tb=12'h0f1;#1; sino_tb=12'h0ee;#1; sino_tb=12'h0eb;#1; sino_tb=12'h0e8;#1; sino_tb=12'h0e5;#1; 
sino_tb=12'h0e2;#1; sino_tb=12'h0df;#1; sino_tb=12'h0db;#1; sino_tb=12'h0d8;#1; sino_tb=12'h0d5;#1; sino_tb=12'h0d2;#1; sino_tb=12'h0cf;#1; sino_tb=12'h0cc;#1; 
sino_tb=12'h0c9;#1; sino_tb=12'h0c6;#1; sino_tb=12'h0c2;#1; sino_tb=12'h0bf;#1; sino_tb=12'h0bc;#1; sino_tb=12'h0b9;#1; sino_tb=12'h0b6;#1; sino_tb=12'h0b3;#1; 
sino_tb=12'h0b0;#1; sino_tb=12'h0ac;#1; sino_tb=12'h0a9;#1; sino_tb=12'h0a6;#1; sino_tb=12'h0a3;#1; sino_tb=12'h0a0;#1; sino_tb=12'h09d;#1; sino_tb=12'h09a;#1; 
sino_tb=12'h097;#1; sino_tb=12'h093;#1; sino_tb=12'h090;#1; sino_tb=12'h08d;#1; sino_tb=12'h08a;#1; sino_tb=12'h087;#1; sino_tb=12'h084;#1; sino_tb=12'h081;#1; 
sino_tb=12'h07e;#1; sino_tb=12'h07a;#1; sino_tb=12'h077;#1; sino_tb=12'h074;#1; sino_tb=12'h071;#1; sino_tb=12'h06e;#1; sino_tb=12'h06b;#1; sino_tb=12'h068;#1; 
sino_tb=12'h064;#1; sino_tb=12'h061;#1; sino_tb=12'h05e;#1; sino_tb=12'h05b;#1; sino_tb=12'h058;#1; sino_tb=12'h055;#1; sino_tb=12'h052;#1; sino_tb=12'h04e;#1; 
sino_tb=12'h04b;#1; sino_tb=12'h048;#1; sino_tb=12'h045;#1; sino_tb=12'h042;#1; sino_tb=12'h03f;#1; sino_tb=12'h03c;#1; sino_tb=12'h039;#1; sino_tb=12'h035;#1; 
sino_tb=12'h032;#1; sino_tb=12'h02f;#1; sino_tb=12'h02c;#1; sino_tb=12'h029;#1; sino_tb=12'h026;#1; sino_tb=12'h023;#1; sino_tb=12'h01f;#1; sino_tb=12'h01c;#1; 
sino_tb=12'h019;#1; sino_tb=12'h016;#1; sino_tb=12'h013;#1; sino_tb=12'h010;#1; sino_tb=12'h00d;#1; sino_tb=12'h009;#1; sino_tb=12'h006;#1; sino_tb=12'h003;#1; 
sino_tb=12'h000;#1; sino_tb=12'hffd;#1; sino_tb=12'hffa;#1; sino_tb=12'hff7;#1; sino_tb=12'hff3;#1; sino_tb=12'hff0;#1; sino_tb=12'hfed;#1; sino_tb=12'hfea;#1; 
sino_tb=12'hfe7;#1; sino_tb=12'hfe4;#1; sino_tb=12'hfe1;#1; sino_tb=12'hfdd;#1; sino_tb=12'hfda;#1; sino_tb=12'hfd7;#1; sino_tb=12'hfd4;#1; sino_tb=12'hfd1;#1; 
sino_tb=12'hfce;#1; sino_tb=12'hfcb;#1; sino_tb=12'hfc7;#1; sino_tb=12'hfc4;#1; sino_tb=12'hfc1;#1; sino_tb=12'hfbe;#1; sino_tb=12'hfbb;#1; sino_tb=12'hfb8;#1; 
sino_tb=12'hfb5;#1; sino_tb=12'hfb2;#1; sino_tb=12'hfae;#1; sino_tb=12'hfab;#1; sino_tb=12'hfa8;#1; sino_tb=12'hfa5;#1; sino_tb=12'hfa2;#1; sino_tb=12'hf9f;#1; 
sino_tb=12'hf9c;#1; sino_tb=12'hf98;#1; sino_tb=12'hf95;#1; sino_tb=12'hf92;#1; sino_tb=12'hf8f;#1; sino_tb=12'hf8c;#1; sino_tb=12'hf89;#1; sino_tb=12'hf86;#1; 
sino_tb=12'hf82;#1; sino_tb=12'hf7f;#1; sino_tb=12'hf7c;#1; sino_tb=12'hf79;#1; sino_tb=12'hf76;#1; sino_tb=12'hf73;#1; sino_tb=12'hf70;#1; sino_tb=12'hf6d;#1; 
sino_tb=12'hf69;#1; sino_tb=12'hf66;#1; sino_tb=12'hf63;#1; sino_tb=12'hf60;#1; sino_tb=12'hf5d;#1; sino_tb=12'hf5a;#1; sino_tb=12'hf57;#1; sino_tb=12'hf54;#1; 
sino_tb=12'hf50;#1; sino_tb=12'hf4d;#1; sino_tb=12'hf4a;#1; sino_tb=12'hf47;#1; sino_tb=12'hf44;#1; sino_tb=12'hf41;#1; sino_tb=12'hf3e;#1; sino_tb=12'hf3a;#1; 
sino_tb=12'hf37;#1; sino_tb=12'hf34;#1; sino_tb=12'hf31;#1; sino_tb=12'hf2e;#1; sino_tb=12'hf2b;#1; sino_tb=12'hf28;#1; sino_tb=12'hf25;#1; sino_tb=12'hf21;#1; 
sino_tb=12'hf1e;#1; sino_tb=12'hf1b;#1; sino_tb=12'hf18;#1; sino_tb=12'hf15;#1; sino_tb=12'hf12;#1; sino_tb=12'hf0f;#1; sino_tb=12'hf0c;#1; sino_tb=12'hf09;#1; 
sino_tb=12'hf05;#1; sino_tb=12'hf02;#1; sino_tb=12'heff;#1; sino_tb=12'hefc;#1; sino_tb=12'hef9;#1; sino_tb=12'hef6;#1; sino_tb=12'hef3;#1; sino_tb=12'hef0;#1; 
sino_tb=12'heed;#1; sino_tb=12'hee9;#1; sino_tb=12'hee6;#1; sino_tb=12'hee3;#1; sino_tb=12'hee0;#1; sino_tb=12'hedd;#1; sino_tb=12'heda;#1; sino_tb=12'hed7;#1; 
sino_tb=12'hed4;#1; sino_tb=12'hed1;#1; sino_tb=12'hecd;#1; sino_tb=12'heca;#1; sino_tb=12'hec7;#1; sino_tb=12'hec4;#1; sino_tb=12'hec1;#1; sino_tb=12'hebe;#1; 
sino_tb=12'hebb;#1; sino_tb=12'heb8;#1; sino_tb=12'heb5;#1; sino_tb=12'heb2;#1; sino_tb=12'heae;#1; sino_tb=12'heab;#1; sino_tb=12'hea8;#1; sino_tb=12'hea5;#1; 
sino_tb=12'hea2;#1; sino_tb=12'he9f;#1; sino_tb=12'he9c;#1; sino_tb=12'he99;#1; sino_tb=12'he96;#1; sino_tb=12'he93;#1; sino_tb=12'he8f;#1; sino_tb=12'he8c;#1; 
sino_tb=12'he89;#1; sino_tb=12'he86;#1; sino_tb=12'he83;#1; sino_tb=12'he80;#1; sino_tb=12'he7d;#1; sino_tb=12'he7a;#1; sino_tb=12'he77;#1; sino_tb=12'he74;#1; 
sino_tb=12'he71;#1; sino_tb=12'he6e;#1; sino_tb=12'he6a;#1; sino_tb=12'he67;#1; sino_tb=12'he64;#1; sino_tb=12'he61;#1; sino_tb=12'he5e;#1; sino_tb=12'he5b;#1; 
sino_tb=12'he58;#1; sino_tb=12'he55;#1; sino_tb=12'he52;#1; sino_tb=12'he4f;#1; sino_tb=12'he4c;#1; sino_tb=12'he49;#1; sino_tb=12'he46;#1; sino_tb=12'he43;#1; 
sino_tb=12'he3f;#1; sino_tb=12'he3c;#1; sino_tb=12'he39;#1; sino_tb=12'he36;#1; sino_tb=12'he33;#1; sino_tb=12'he30;#1; sino_tb=12'he2d;#1; sino_tb=12'he2a;#1; 
sino_tb=12'he27;#1; sino_tb=12'he24;#1; sino_tb=12'he21;#1; sino_tb=12'he1e;#1; sino_tb=12'he1b;#1; sino_tb=12'he18;#1; sino_tb=12'he15;#1; sino_tb=12'he12;#1; 
sino_tb=12'he0f;#1; sino_tb=12'he0c;#1; sino_tb=12'he09;#1; sino_tb=12'he05;#1; sino_tb=12'he02;#1; sino_tb=12'hdff;#1; sino_tb=12'hdfc;#1; sino_tb=12'hdf9;#1; 
sino_tb=12'hdf6;#1; sino_tb=12'hdf3;#1; sino_tb=12'hdf0;#1; sino_tb=12'hded;#1; sino_tb=12'hdea;#1; sino_tb=12'hde7;#1; sino_tb=12'hde4;#1; sino_tb=12'hde1;#1; 
sino_tb=12'hdde;#1; sino_tb=12'hddb;#1; sino_tb=12'hdd8;#1; sino_tb=12'hdd5;#1; sino_tb=12'hdd2;#1; sino_tb=12'hdcf;#1; sino_tb=12'hdcc;#1; sino_tb=12'hdc9;#1; 
sino_tb=12'hdc6;#1; sino_tb=12'hdc3;#1; sino_tb=12'hdc0;#1; sino_tb=12'hdbd;#1; sino_tb=12'hdba;#1; sino_tb=12'hdb7;#1; sino_tb=12'hdb4;#1; sino_tb=12'hdb1;#1; 
sino_tb=12'hdae;#1; sino_tb=12'hdab;#1; sino_tb=12'hda8;#1; sino_tb=12'hda5;#1; sino_tb=12'hda2;#1; sino_tb=12'hd9f;#1; sino_tb=12'hd9c;#1; sino_tb=12'hd99;#1; 
sino_tb=12'hd96;#1; sino_tb=12'hd93;#1; sino_tb=12'hd90;#1; sino_tb=12'hd8d;#1; sino_tb=12'hd8a;#1; sino_tb=12'hd87;#1; sino_tb=12'hd84;#1; sino_tb=12'hd81;#1; 
sino_tb=12'hd7e;#1; sino_tb=12'hd7b;#1; sino_tb=12'hd78;#1; sino_tb=12'hd75;#1; sino_tb=12'hd72;#1; sino_tb=12'hd6f;#1; sino_tb=12'hd6c;#1; sino_tb=12'hd69;#1; 
sino_tb=12'hd66;#1; sino_tb=12'hd63;#1; sino_tb=12'hd60;#1; sino_tb=12'hd5d;#1; sino_tb=12'hd5a;#1; sino_tb=12'hd57;#1; sino_tb=12'hd54;#1; sino_tb=12'hd51;#1; 
sino_tb=12'hd4e;#1; sino_tb=12'hd4b;#1; sino_tb=12'hd48;#1; sino_tb=12'hd46;#1; sino_tb=12'hd43;#1; sino_tb=12'hd40;#1; sino_tb=12'hd3d;#1; sino_tb=12'hd3a;#1; 
sino_tb=12'hd37;#1; sino_tb=12'hd34;#1; sino_tb=12'hd31;#1; sino_tb=12'hd2e;#1; sino_tb=12'hd2b;#1; sino_tb=12'hd28;#1; sino_tb=12'hd25;#1; sino_tb=12'hd22;#1; 
sino_tb=12'hd1f;#1; sino_tb=12'hd1c;#1; sino_tb=12'hd19;#1; sino_tb=12'hd17;#1; sino_tb=12'hd14;#1; sino_tb=12'hd11;#1; sino_tb=12'hd0e;#1; sino_tb=12'hd0b;#1; 
sino_tb=12'hd08;#1; sino_tb=12'hd05;#1; sino_tb=12'hd02;#1; sino_tb=12'hcff;#1; sino_tb=12'hcfc;#1; sino_tb=12'hcf9;#1; sino_tb=12'hcf6;#1; sino_tb=12'hcf4;#1; 
sino_tb=12'hcf1;#1; sino_tb=12'hcee;#1; sino_tb=12'hceb;#1; sino_tb=12'hce8;#1; sino_tb=12'hce5;#1; sino_tb=12'hce2;#1; sino_tb=12'hcdf;#1; sino_tb=12'hcdc;#1; 
sino_tb=12'hcd9;#1; sino_tb=12'hcd7;#1; sino_tb=12'hcd4;#1; sino_tb=12'hcd1;#1; sino_tb=12'hcce;#1; sino_tb=12'hccb;#1; sino_tb=12'hcc8;#1; sino_tb=12'hcc5;#1; 
sino_tb=12'hcc2;#1; sino_tb=12'hcc0;#1; sino_tb=12'hcbd;#1; sino_tb=12'hcba;#1; sino_tb=12'hcb7;#1; sino_tb=12'hcb4;#1; sino_tb=12'hcb1;#1; sino_tb=12'hcae;#1; 
sino_tb=12'hcac;#1; sino_tb=12'hca9;#1; sino_tb=12'hca6;#1; sino_tb=12'hca3;#1; sino_tb=12'hca0;#1; sino_tb=12'hc9d;#1; sino_tb=12'hc9a;#1; sino_tb=12'hc98;#1; 
sino_tb=12'hc95;#1; sino_tb=12'hc92;#1; sino_tb=12'hc8f;#1; sino_tb=12'hc8c;#1; sino_tb=12'hc89;#1; sino_tb=12'hc87;#1; sino_tb=12'hc84;#1; sino_tb=12'hc81;#1; 
sino_tb=12'hc7e;#1; sino_tb=12'hc7b;#1; sino_tb=12'hc79;#1; sino_tb=12'hc76;#1; sino_tb=12'hc73;#1; sino_tb=12'hc70;#1; sino_tb=12'hc6d;#1; sino_tb=12'hc6a;#1; 
sino_tb=12'hc68;#1; sino_tb=12'hc65;#1; sino_tb=12'hc62;#1; sino_tb=12'hc5f;#1; sino_tb=12'hc5c;#1; sino_tb=12'hc5a;#1; sino_tb=12'hc57;#1; sino_tb=12'hc54;#1; 
sino_tb=12'hc51;#1; sino_tb=12'hc4e;#1; sino_tb=12'hc4c;#1; sino_tb=12'hc49;#1; sino_tb=12'hc46;#1; sino_tb=12'hc43;#1; sino_tb=12'hc41;#1; sino_tb=12'hc3e;#1; 
sino_tb=12'hc3b;#1; sino_tb=12'hc38;#1; sino_tb=12'hc36;#1; sino_tb=12'hc33;#1; sino_tb=12'hc30;#1; sino_tb=12'hc2d;#1; sino_tb=12'hc2a;#1; sino_tb=12'hc28;#1; 
sino_tb=12'hc25;#1; sino_tb=12'hc22;#1; sino_tb=12'hc1f;#1; sino_tb=12'hc1d;#1; sino_tb=12'hc1a;#1; sino_tb=12'hc17;#1; sino_tb=12'hc15;#1; sino_tb=12'hc12;#1; 
sino_tb=12'hc0f;#1; sino_tb=12'hc0c;#1; sino_tb=12'hc0a;#1; sino_tb=12'hc07;#1; sino_tb=12'hc04;#1; sino_tb=12'hc01;#1; sino_tb=12'hbff;#1; sino_tb=12'hbfc;#1; 
sino_tb=12'hbf9;#1; sino_tb=12'hbf7;#1; sino_tb=12'hbf4;#1; sino_tb=12'hbf1;#1; sino_tb=12'hbee;#1; sino_tb=12'hbec;#1; sino_tb=12'hbe9;#1; sino_tb=12'hbe6;#1; 
sino_tb=12'hbe4;#1; sino_tb=12'hbe1;#1; sino_tb=12'hbde;#1; sino_tb=12'hbdc;#1; sino_tb=12'hbd9;#1; sino_tb=12'hbd6;#1; sino_tb=12'hbd4;#1; sino_tb=12'hbd1;#1; 
sino_tb=12'hbce;#1; sino_tb=12'hbcb;#1; sino_tb=12'hbc9;#1; sino_tb=12'hbc6;#1; sino_tb=12'hbc3;#1; sino_tb=12'hbc1;#1; sino_tb=12'hbbe;#1; sino_tb=12'hbbc;#1; 
sino_tb=12'hbb9;#1; sino_tb=12'hbb6;#1; sino_tb=12'hbb4;#1; sino_tb=12'hbb1;#1; sino_tb=12'hbae;#1; sino_tb=12'hbac;#1; sino_tb=12'hba9;#1; sino_tb=12'hba6;#1; 
sino_tb=12'hba4;#1; sino_tb=12'hba1;#1; sino_tb=12'hb9e;#1; sino_tb=12'hb9c;#1; sino_tb=12'hb99;#1; sino_tb=12'hb97;#1; sino_tb=12'hb94;#1; sino_tb=12'hb91;#1; 
sino_tb=12'hb8f;#1; sino_tb=12'hb8c;#1; sino_tb=12'hb8a;#1; sino_tb=12'hb87;#1; sino_tb=12'hb84;#1; sino_tb=12'hb82;#1; sino_tb=12'hb7f;#1; sino_tb=12'hb7d;#1; 
sino_tb=12'hb7a;#1; sino_tb=12'hb77;#1; sino_tb=12'hb75;#1; sino_tb=12'hb72;#1; sino_tb=12'hb70;#1; sino_tb=12'hb6d;#1; sino_tb=12'hb6a;#1; sino_tb=12'hb68;#1; 
sino_tb=12'hb65;#1; sino_tb=12'hb63;#1; sino_tb=12'hb60;#1; sino_tb=12'hb5e;#1; sino_tb=12'hb5b;#1; sino_tb=12'hb59;#1; sino_tb=12'hb56;#1; sino_tb=12'hb53;#1; 
sino_tb=12'hb51;#1; sino_tb=12'hb4e;#1; sino_tb=12'hb4c;#1; sino_tb=12'hb49;#1; sino_tb=12'hb47;#1; sino_tb=12'hb44;#1; sino_tb=12'hb42;#1; sino_tb=12'hb3f;#1; 
sino_tb=12'hb3d;#1; sino_tb=12'hb3a;#1; sino_tb=12'hb38;#1; sino_tb=12'hb35;#1; sino_tb=12'hb33;#1; sino_tb=12'hb30;#1; sino_tb=12'hb2e;#1; sino_tb=12'hb2b;#1; 
sino_tb=12'hb29;#1; sino_tb=12'hb26;#1; sino_tb=12'hb24;#1; sino_tb=12'hb21;#1; sino_tb=12'hb1f;#1; sino_tb=12'hb1c;#1; sino_tb=12'hb1a;#1; sino_tb=12'hb17;#1; 
sino_tb=12'hb15;#1; sino_tb=12'hb12;#1; sino_tb=12'hb10;#1; sino_tb=12'hb0d;#1; sino_tb=12'hb0b;#1; sino_tb=12'hb08;#1; sino_tb=12'hb06;#1; sino_tb=12'hb03;#1; 
sino_tb=12'hb01;#1; sino_tb=12'hafe;#1; sino_tb=12'hafc;#1; sino_tb=12'hafa;#1; sino_tb=12'haf7;#1; sino_tb=12'haf5;#1; sino_tb=12'haf2;#1; sino_tb=12'haf0;#1; 
sino_tb=12'haed;#1; sino_tb=12'haeb;#1; sino_tb=12'hae9;#1; sino_tb=12'hae6;#1; sino_tb=12'hae4;#1; sino_tb=12'hae1;#1; sino_tb=12'hadf;#1; sino_tb=12'hadc;#1; 
sino_tb=12'hada;#1; sino_tb=12'had8;#1; sino_tb=12'had5;#1; sino_tb=12'had3;#1; sino_tb=12'had0;#1; sino_tb=12'hace;#1; sino_tb=12'hacc;#1; sino_tb=12'hac9;#1; 
sino_tb=12'hac7;#1; sino_tb=12'hac5;#1; sino_tb=12'hac2;#1; sino_tb=12'hac0;#1; sino_tb=12'habd;#1; sino_tb=12'habb;#1; sino_tb=12'hab9;#1; sino_tb=12'hab6;#1; 
sino_tb=12'hab4;#1; sino_tb=12'hab2;#1; sino_tb=12'haaf;#1; sino_tb=12'haad;#1; sino_tb=12'haab;#1; sino_tb=12'haa8;#1; sino_tb=12'haa6;#1; sino_tb=12'haa4;#1; 
sino_tb=12'haa1;#1; sino_tb=12'ha9f;#1; sino_tb=12'ha9d;#1; sino_tb=12'ha9a;#1; sino_tb=12'ha98;#1; sino_tb=12'ha96;#1; sino_tb=12'ha93;#1; sino_tb=12'ha91;#1; 
sino_tb=12'ha8f;#1; sino_tb=12'ha8d;#1; sino_tb=12'ha8a;#1; sino_tb=12'ha88;#1; sino_tb=12'ha86;#1; sino_tb=12'ha83;#1; sino_tb=12'ha81;#1; sino_tb=12'ha7f;#1; 
sino_tb=12'ha7d;#1; sino_tb=12'ha7a;#1; sino_tb=12'ha78;#1; sino_tb=12'ha76;#1; sino_tb=12'ha73;#1; sino_tb=12'ha71;#1; sino_tb=12'ha6f;#1; sino_tb=12'ha6d;#1; 
sino_tb=12'ha6a;#1; sino_tb=12'ha68;#1; sino_tb=12'ha66;#1; sino_tb=12'ha64;#1; sino_tb=12'ha61;#1; sino_tb=12'ha5f;#1; sino_tb=12'ha5d;#1; sino_tb=12'ha5b;#1; 
sino_tb=12'ha59;#1; sino_tb=12'ha56;#1; sino_tb=12'ha54;#1; sino_tb=12'ha52;#1; sino_tb=12'ha50;#1; sino_tb=12'ha4d;#1; sino_tb=12'ha4b;#1; sino_tb=12'ha49;#1; 
sino_tb=12'ha47;#1; sino_tb=12'ha45;#1; sino_tb=12'ha43;#1; sino_tb=12'ha40;#1; sino_tb=12'ha3e;#1; sino_tb=12'ha3c;#1; sino_tb=12'ha3a;#1; sino_tb=12'ha38;#1; 
sino_tb=12'ha35;#1; sino_tb=12'ha33;#1; sino_tb=12'ha31;#1; sino_tb=12'ha2f;#1; sino_tb=12'ha2d;#1; sino_tb=12'ha2b;#1; sino_tb=12'ha29;#1; sino_tb=12'ha26;#1; 
sino_tb=12'ha24;#1; sino_tb=12'ha22;#1; sino_tb=12'ha20;#1; sino_tb=12'ha1e;#1; sino_tb=12'ha1c;#1; sino_tb=12'ha1a;#1; sino_tb=12'ha17;#1; sino_tb=12'ha15;#1; 
sino_tb=12'ha13;#1; sino_tb=12'ha11;#1; sino_tb=12'ha0f;#1; sino_tb=12'ha0d;#1; sino_tb=12'ha0b;#1; sino_tb=12'ha09;#1; sino_tb=12'ha07;#1; sino_tb=12'ha05;#1; 
sino_tb=12'ha03;#1; sino_tb=12'ha00;#1; sino_tb=12'h9fe;#1; sino_tb=12'h9fc;#1; sino_tb=12'h9fa;#1; sino_tb=12'h9f8;#1; sino_tb=12'h9f6;#1; sino_tb=12'h9f4;#1; 
sino_tb=12'h9f2;#1; sino_tb=12'h9f0;#1; sino_tb=12'h9ee;#1; sino_tb=12'h9ec;#1; sino_tb=12'h9ea;#1; sino_tb=12'h9e8;#1; sino_tb=12'h9e6;#1; sino_tb=12'h9e4;#1; 
sino_tb=12'h9e2;#1; sino_tb=12'h9e0;#1; sino_tb=12'h9de;#1; sino_tb=12'h9dc;#1; sino_tb=12'h9da;#1; sino_tb=12'h9d8;#1; sino_tb=12'h9d6;#1; sino_tb=12'h9d4;#1; 
sino_tb=12'h9d2;#1; sino_tb=12'h9d0;#1; sino_tb=12'h9ce;#1; sino_tb=12'h9cc;#1; sino_tb=12'h9ca;#1; sino_tb=12'h9c8;#1; sino_tb=12'h9c6;#1; sino_tb=12'h9c4;#1; 
sino_tb=12'h9c2;#1; sino_tb=12'h9c0;#1; sino_tb=12'h9be;#1; sino_tb=12'h9bc;#1; sino_tb=12'h9ba;#1; sino_tb=12'h9b8;#1; sino_tb=12'h9b6;#1; sino_tb=12'h9b4;#1; 
sino_tb=12'h9b2;#1; sino_tb=12'h9b0;#1; sino_tb=12'h9ae;#1; sino_tb=12'h9ac;#1; sino_tb=12'h9ab;#1; sino_tb=12'h9a9;#1; sino_tb=12'h9a7;#1; sino_tb=12'h9a5;#1; 
sino_tb=12'h9a3;#1; sino_tb=12'h9a1;#1; sino_tb=12'h99f;#1; sino_tb=12'h99d;#1; sino_tb=12'h99b;#1; sino_tb=12'h999;#1; sino_tb=12'h998;#1; sino_tb=12'h996;#1; 
sino_tb=12'h994;#1; sino_tb=12'h992;#1; sino_tb=12'h990;#1; sino_tb=12'h98e;#1; sino_tb=12'h98c;#1; sino_tb=12'h98b;#1; sino_tb=12'h989;#1; sino_tb=12'h987;#1; 
sino_tb=12'h985;#1; sino_tb=12'h983;#1; sino_tb=12'h981;#1; sino_tb=12'h97f;#1; sino_tb=12'h97e;#1; sino_tb=12'h97c;#1; sino_tb=12'h97a;#1; sino_tb=12'h978;#1; 
sino_tb=12'h976;#1; sino_tb=12'h975;#1; sino_tb=12'h973;#1; sino_tb=12'h971;#1; sino_tb=12'h96f;#1; sino_tb=12'h96d;#1; sino_tb=12'h96c;#1; sino_tb=12'h96a;#1; 
sino_tb=12'h968;#1; sino_tb=12'h966;#1; sino_tb=12'h965;#1; sino_tb=12'h963;#1; sino_tb=12'h961;#1; sino_tb=12'h95f;#1; sino_tb=12'h95d;#1; sino_tb=12'h95c;#1; 
sino_tb=12'h95a;#1; sino_tb=12'h958;#1; sino_tb=12'h957;#1; sino_tb=12'h955;#1; sino_tb=12'h953;#1; sino_tb=12'h951;#1; sino_tb=12'h950;#1; sino_tb=12'h94e;#1; 
sino_tb=12'h94c;#1; sino_tb=12'h94a;#1; sino_tb=12'h949;#1; sino_tb=12'h947;#1; sino_tb=12'h945;#1; sino_tb=12'h944;#1; sino_tb=12'h942;#1; sino_tb=12'h940;#1; 
sino_tb=12'h93f;#1; sino_tb=12'h93d;#1; sino_tb=12'h93b;#1; sino_tb=12'h93a;#1; sino_tb=12'h938;#1; sino_tb=12'h936;#1; sino_tb=12'h935;#1; sino_tb=12'h933;#1; 
sino_tb=12'h931;#1; sino_tb=12'h930;#1; sino_tb=12'h92e;#1; sino_tb=12'h92c;#1; sino_tb=12'h92b;#1; sino_tb=12'h929;#1; sino_tb=12'h927;#1; sino_tb=12'h926;#1; 
sino_tb=12'h924;#1; sino_tb=12'h923;#1; sino_tb=12'h921;#1; sino_tb=12'h91f;#1; sino_tb=12'h91e;#1; sino_tb=12'h91c;#1; sino_tb=12'h91b;#1; sino_tb=12'h919;#1; 
sino_tb=12'h917;#1; sino_tb=12'h916;#1; sino_tb=12'h914;#1; sino_tb=12'h913;#1; sino_tb=12'h911;#1; sino_tb=12'h910;#1; sino_tb=12'h90e;#1; sino_tb=12'h90c;#1; 
sino_tb=12'h90b;#1; sino_tb=12'h909;#1; sino_tb=12'h908;#1; sino_tb=12'h906;#1; sino_tb=12'h905;#1; sino_tb=12'h903;#1; sino_tb=12'h902;#1; sino_tb=12'h900;#1; 
sino_tb=12'h8ff;#1; sino_tb=12'h8fd;#1; sino_tb=12'h8fc;#1; sino_tb=12'h8fa;#1; sino_tb=12'h8f9;#1; sino_tb=12'h8f7;#1; sino_tb=12'h8f6;#1; sino_tb=12'h8f4;#1; 
sino_tb=12'h8f3;#1; sino_tb=12'h8f1;#1; sino_tb=12'h8f0;#1; sino_tb=12'h8ee;#1; sino_tb=12'h8ed;#1; sino_tb=12'h8eb;#1; sino_tb=12'h8ea;#1; sino_tb=12'h8e8;#1; 
sino_tb=12'h8e7;#1; sino_tb=12'h8e6;#1; sino_tb=12'h8e4;#1; sino_tb=12'h8e3;#1; sino_tb=12'h8e1;#1; sino_tb=12'h8e0;#1; sino_tb=12'h8de;#1; sino_tb=12'h8dd;#1; 
sino_tb=12'h8dc;#1; sino_tb=12'h8da;#1; sino_tb=12'h8d9;#1; sino_tb=12'h8d7;#1; sino_tb=12'h8d6;#1; sino_tb=12'h8d5;#1; sino_tb=12'h8d3;#1; sino_tb=12'h8d2;#1; 
sino_tb=12'h8d0;#1; sino_tb=12'h8cf;#1; sino_tb=12'h8ce;#1; sino_tb=12'h8cc;#1; sino_tb=12'h8cb;#1; sino_tb=12'h8ca;#1; sino_tb=12'h8c8;#1; sino_tb=12'h8c7;#1; 
sino_tb=12'h8c6;#1; sino_tb=12'h8c4;#1; sino_tb=12'h8c3;#1; sino_tb=12'h8c2;#1; sino_tb=12'h8c0;#1; sino_tb=12'h8bf;#1; sino_tb=12'h8be;#1; sino_tb=12'h8bc;#1; 
sino_tb=12'h8bb;#1; sino_tb=12'h8ba;#1; sino_tb=12'h8b8;#1; sino_tb=12'h8b7;#1; sino_tb=12'h8b6;#1; sino_tb=12'h8b4;#1; sino_tb=12'h8b3;#1; sino_tb=12'h8b2;#1; 
sino_tb=12'h8b1;#1; sino_tb=12'h8af;#1; sino_tb=12'h8ae;#1; sino_tb=12'h8ad;#1; sino_tb=12'h8ac;#1; sino_tb=12'h8aa;#1; sino_tb=12'h8a9;#1; sino_tb=12'h8a8;#1; 
sino_tb=12'h8a7;#1; sino_tb=12'h8a5;#1; sino_tb=12'h8a4;#1; sino_tb=12'h8a3;#1; sino_tb=12'h8a2;#1; sino_tb=12'h8a0;#1; sino_tb=12'h89f;#1; sino_tb=12'h89e;#1; 
sino_tb=12'h89d;#1; sino_tb=12'h89c;#1; sino_tb=12'h89a;#1; sino_tb=12'h899;#1; sino_tb=12'h898;#1; sino_tb=12'h897;#1; sino_tb=12'h896;#1; sino_tb=12'h895;#1; 
sino_tb=12'h893;#1; sino_tb=12'h892;#1; sino_tb=12'h891;#1; sino_tb=12'h890;#1; sino_tb=12'h88f;#1; sino_tb=12'h88e;#1; sino_tb=12'h88c;#1; sino_tb=12'h88b;#1; 
sino_tb=12'h88a;#1; sino_tb=12'h889;#1; sino_tb=12'h888;#1; sino_tb=12'h887;#1; sino_tb=12'h886;#1; sino_tb=12'h885;#1; sino_tb=12'h883;#1; sino_tb=12'h882;#1; 
sino_tb=12'h881;#1; sino_tb=12'h880;#1; sino_tb=12'h87f;#1; sino_tb=12'h87e;#1; sino_tb=12'h87d;#1; sino_tb=12'h87c;#1; sino_tb=12'h87b;#1; sino_tb=12'h87a;#1; 
sino_tb=12'h879;#1; sino_tb=12'h878;#1; sino_tb=12'h877;#1; sino_tb=12'h876;#1; sino_tb=12'h874;#1; sino_tb=12'h873;#1; sino_tb=12'h872;#1; sino_tb=12'h871;#1; 
sino_tb=12'h870;#1; sino_tb=12'h86f;#1; sino_tb=12'h86e;#1; sino_tb=12'h86d;#1; sino_tb=12'h86c;#1; sino_tb=12'h86b;#1; sino_tb=12'h86a;#1; sino_tb=12'h869;#1; 
sino_tb=12'h868;#1; sino_tb=12'h867;#1; sino_tb=12'h866;#1; sino_tb=12'h865;#1; sino_tb=12'h864;#1; sino_tb=12'h863;#1; sino_tb=12'h862;#1; sino_tb=12'h862;#1; 
sino_tb=12'h861;#1; sino_tb=12'h860;#1; sino_tb=12'h85f;#1; sino_tb=12'h85e;#1; sino_tb=12'h85d;#1; sino_tb=12'h85c;#1; sino_tb=12'h85b;#1; sino_tb=12'h85a;#1; 
sino_tb=12'h859;#1; sino_tb=12'h858;#1; sino_tb=12'h857;#1; sino_tb=12'h856;#1; sino_tb=12'h856;#1; sino_tb=12'h855;#1; sino_tb=12'h854;#1; sino_tb=12'h853;#1; 
sino_tb=12'h852;#1; sino_tb=12'h851;#1; sino_tb=12'h850;#1; sino_tb=12'h84f;#1; sino_tb=12'h84f;#1; sino_tb=12'h84e;#1; sino_tb=12'h84d;#1; sino_tb=12'h84c;#1; 
sino_tb=12'h84b;#1; sino_tb=12'h84a;#1; sino_tb=12'h849;#1; sino_tb=12'h849;#1; sino_tb=12'h848;#1; sino_tb=12'h847;#1; sino_tb=12'h846;#1; sino_tb=12'h845;#1; 
sino_tb=12'h845;#1; sino_tb=12'h844;#1; sino_tb=12'h843;#1; sino_tb=12'h842;#1; sino_tb=12'h841;#1; sino_tb=12'h841;#1; sino_tb=12'h840;#1; sino_tb=12'h83f;#1; 
sino_tb=12'h83e;#1; sino_tb=12'h83e;#1; sino_tb=12'h83d;#1; sino_tb=12'h83c;#1; sino_tb=12'h83b;#1; sino_tb=12'h83b;#1; sino_tb=12'h83a;#1; sino_tb=12'h839;#1; 
sino_tb=12'h838;#1; sino_tb=12'h838;#1; sino_tb=12'h837;#1; sino_tb=12'h836;#1; sino_tb=12'h836;#1; sino_tb=12'h835;#1; sino_tb=12'h834;#1; sino_tb=12'h833;#1; 
sino_tb=12'h833;#1; sino_tb=12'h832;#1; sino_tb=12'h831;#1; sino_tb=12'h831;#1; sino_tb=12'h830;#1; sino_tb=12'h82f;#1; sino_tb=12'h82f;#1; sino_tb=12'h82e;#1; 
sino_tb=12'h82d;#1; sino_tb=12'h82d;#1; sino_tb=12'h82c;#1; sino_tb=12'h82b;#1; sino_tb=12'h82b;#1; sino_tb=12'h82a;#1; sino_tb=12'h82a;#1; sino_tb=12'h829;#1; 
sino_tb=12'h828;#1; sino_tb=12'h828;#1; sino_tb=12'h827;#1; sino_tb=12'h827;#1; sino_tb=12'h826;#1; sino_tb=12'h825;#1; sino_tb=12'h825;#1; sino_tb=12'h824;#1; 
sino_tb=12'h824;#1; sino_tb=12'h823;#1; sino_tb=12'h822;#1; sino_tb=12'h822;#1; sino_tb=12'h821;#1; sino_tb=12'h821;#1; sino_tb=12'h820;#1; sino_tb=12'h820;#1; 
sino_tb=12'h81f;#1; sino_tb=12'h81f;#1; sino_tb=12'h81e;#1; sino_tb=12'h81e;#1; sino_tb=12'h81d;#1; sino_tb=12'h81d;#1; sino_tb=12'h81c;#1; sino_tb=12'h81b;#1; 
sino_tb=12'h81b;#1; sino_tb=12'h81a;#1; sino_tb=12'h81a;#1; sino_tb=12'h81a;#1; sino_tb=12'h819;#1; sino_tb=12'h819;#1; sino_tb=12'h818;#1; sino_tb=12'h818;#1; 
sino_tb=12'h817;#1; sino_tb=12'h817;#1; sino_tb=12'h816;#1; sino_tb=12'h816;#1; sino_tb=12'h815;#1; sino_tb=12'h815;#1; sino_tb=12'h814;#1; sino_tb=12'h814;#1; 
sino_tb=12'h814;#1; sino_tb=12'h813;#1; sino_tb=12'h813;#1; sino_tb=12'h812;#1; sino_tb=12'h812;#1; sino_tb=12'h812;#1; sino_tb=12'h811;#1; sino_tb=12'h811;#1; 
sino_tb=12'h810;#1; sino_tb=12'h810;#1; sino_tb=12'h810;#1; sino_tb=12'h80f;#1; sino_tb=12'h80f;#1; sino_tb=12'h80f;#1; sino_tb=12'h80e;#1; sino_tb=12'h80e;#1; 
sino_tb=12'h80d;#1; sino_tb=12'h80d;#1; sino_tb=12'h80d;#1; sino_tb=12'h80c;#1; sino_tb=12'h80c;#1; sino_tb=12'h80c;#1; sino_tb=12'h80b;#1; sino_tb=12'h80b;#1; 
sino_tb=12'h80b;#1; sino_tb=12'h80b;#1; sino_tb=12'h80a;#1; sino_tb=12'h80a;#1; sino_tb=12'h80a;#1; sino_tb=12'h809;#1; sino_tb=12'h809;#1; sino_tb=12'h809;#1; 
sino_tb=12'h809;#1; sino_tb=12'h808;#1; sino_tb=12'h808;#1; sino_tb=12'h808;#1; sino_tb=12'h808;#1; sino_tb=12'h807;#1; sino_tb=12'h807;#1; sino_tb=12'h807;#1; 
sino_tb=12'h807;#1; sino_tb=12'h806;#1; sino_tb=12'h806;#1; sino_tb=12'h806;#1; sino_tb=12'h806;#1; sino_tb=12'h805;#1; sino_tb=12'h805;#1; sino_tb=12'h805;#1; 
sino_tb=12'h805;#1; sino_tb=12'h805;#1; sino_tb=12'h804;#1; sino_tb=12'h804;#1; sino_tb=12'h804;#1; sino_tb=12'h804;#1; sino_tb=12'h804;#1; sino_tb=12'h804;#1; 
sino_tb=12'h803;#1; sino_tb=12'h803;#1; sino_tb=12'h803;#1; sino_tb=12'h803;#1; sino_tb=12'h803;#1; sino_tb=12'h803;#1; sino_tb=12'h803;#1; sino_tb=12'h803;#1; 
sino_tb=12'h802;#1; sino_tb=12'h802;#1; sino_tb=12'h802;#1; sino_tb=12'h802;#1; sino_tb=12'h802;#1; sino_tb=12'h802;#1; sino_tb=12'h802;#1; sino_tb=12'h802;#1; 
sino_tb=12'h802;#1; sino_tb=12'h802;#1; sino_tb=12'h801;#1; sino_tb=12'h801;#1; sino_tb=12'h801;#1; sino_tb=12'h801;#1; sino_tb=12'h801;#1; sino_tb=12'h801;#1; 
sino_tb=12'h801;#1; sino_tb=12'h801;#1; sino_tb=12'h801;#1; sino_tb=12'h801;#1; sino_tb=12'h801;#1; sino_tb=12'h801;#1; sino_tb=12'h801;#1; sino_tb=12'h801;#1; 
sino_tb=12'h801;#1; sino_tb=12'h801;#1; sino_tb=12'h801;#1; sino_tb=12'h801;#1; sino_tb=12'h801;#1; sino_tb=12'h801;#1; sino_tb=12'h801;#1; sino_tb=12'h801;#1; 
sino_tb=12'h801;#1; sino_tb=12'h801;#1; sino_tb=12'h801;#1; sino_tb=12'h801;#1; sino_tb=12'h801;#1; sino_tb=12'h801;#1; sino_tb=12'h801;#1; sino_tb=12'h802;#1; 
sino_tb=12'h802;#1; sino_tb=12'h802;#1; sino_tb=12'h802;#1; sino_tb=12'h802;#1; sino_tb=12'h802;#1; sino_tb=12'h802;#1; sino_tb=12'h802;#1; sino_tb=12'h802;#1; 
sino_tb=12'h802;#1; sino_tb=12'h803;#1; sino_tb=12'h803;#1; sino_tb=12'h803;#1; sino_tb=12'h803;#1; sino_tb=12'h803;#1; sino_tb=12'h803;#1; sino_tb=12'h803;#1; 
sino_tb=12'h803;#1; sino_tb=12'h804;#1; sino_tb=12'h804;#1; sino_tb=12'h804;#1; sino_tb=12'h804;#1; sino_tb=12'h804;#1; sino_tb=12'h804;#1; sino_tb=12'h805;#1; 
sino_tb=12'h805;#1; sino_tb=12'h805;#1; sino_tb=12'h805;#1; sino_tb=12'h805;#1; sino_tb=12'h806;#1; sino_tb=12'h806;#1; sino_tb=12'h806;#1; sino_tb=12'h806;#1; 
sino_tb=12'h807;#1; sino_tb=12'h807;#1; sino_tb=12'h807;#1; sino_tb=12'h807;#1; sino_tb=12'h808;#1; sino_tb=12'h808;#1; sino_tb=12'h808;#1; sino_tb=12'h808;#1; 
sino_tb=12'h809;#1; sino_tb=12'h809;#1; sino_tb=12'h809;#1; sino_tb=12'h809;#1; sino_tb=12'h80a;#1; sino_tb=12'h80a;#1; sino_tb=12'h80a;#1; sino_tb=12'h80b;#1; 
sino_tb=12'h80b;#1; sino_tb=12'h80b;#1; sino_tb=12'h80b;#1; sino_tb=12'h80c;#1; sino_tb=12'h80c;#1; sino_tb=12'h80c;#1; sino_tb=12'h80d;#1; sino_tb=12'h80d;#1; 
sino_tb=12'h80d;#1; sino_tb=12'h80e;#1; sino_tb=12'h80e;#1; sino_tb=12'h80f;#1; sino_tb=12'h80f;#1; sino_tb=12'h80f;#1; sino_tb=12'h810;#1; sino_tb=12'h810;#1; 
sino_tb=12'h810;#1; sino_tb=12'h811;#1; sino_tb=12'h811;#1; sino_tb=12'h812;#1; sino_tb=12'h812;#1; sino_tb=12'h812;#1; sino_tb=12'h813;#1; sino_tb=12'h813;#1; 
sino_tb=12'h814;#1; sino_tb=12'h814;#1; sino_tb=12'h814;#1; sino_tb=12'h815;#1; sino_tb=12'h815;#1; sino_tb=12'h816;#1; sino_tb=12'h816;#1; sino_tb=12'h817;#1; 
sino_tb=12'h817;#1; sino_tb=12'h818;#1; sino_tb=12'h818;#1; sino_tb=12'h819;#1; sino_tb=12'h819;#1; sino_tb=12'h81a;#1; sino_tb=12'h81a;#1; sino_tb=12'h81a;#1; 
sino_tb=12'h81b;#1; sino_tb=12'h81b;#1; sino_tb=12'h81c;#1; sino_tb=12'h81d;#1; sino_tb=12'h81d;#1; sino_tb=12'h81e;#1; sino_tb=12'h81e;#1; sino_tb=12'h81f;#1; 
sino_tb=12'h81f;#1; sino_tb=12'h820;#1; sino_tb=12'h820;#1; sino_tb=12'h821;#1; sino_tb=12'h821;#1; sino_tb=12'h822;#1; sino_tb=12'h822;#1; sino_tb=12'h823;#1; 
sino_tb=12'h824;#1; sino_tb=12'h824;#1; sino_tb=12'h825;#1; sino_tb=12'h825;#1; sino_tb=12'h826;#1; sino_tb=12'h827;#1; sino_tb=12'h827;#1; sino_tb=12'h828;#1; 
sino_tb=12'h828;#1; sino_tb=12'h829;#1; sino_tb=12'h82a;#1; sino_tb=12'h82a;#1; sino_tb=12'h82b;#1; sino_tb=12'h82b;#1; sino_tb=12'h82c;#1; sino_tb=12'h82d;#1; 
sino_tb=12'h82d;#1; sino_tb=12'h82e;#1; sino_tb=12'h82f;#1; sino_tb=12'h82f;#1; sino_tb=12'h830;#1; sino_tb=12'h831;#1; sino_tb=12'h831;#1; sino_tb=12'h832;#1; 
sino_tb=12'h833;#1; sino_tb=12'h833;#1; sino_tb=12'h834;#1; sino_tb=12'h835;#1; sino_tb=12'h836;#1; sino_tb=12'h836;#1; sino_tb=12'h837;#1; sino_tb=12'h838;#1; 
sino_tb=12'h838;#1; sino_tb=12'h839;#1; sino_tb=12'h83a;#1; sino_tb=12'h83b;#1; sino_tb=12'h83b;#1; sino_tb=12'h83c;#1; sino_tb=12'h83d;#1; sino_tb=12'h83e;#1; 
sino_tb=12'h83e;#1; sino_tb=12'h83f;#1; sino_tb=12'h840;#1; sino_tb=12'h841;#1; sino_tb=12'h841;#1; sino_tb=12'h842;#1; sino_tb=12'h843;#1; sino_tb=12'h844;#1; 
sino_tb=12'h845;#1; sino_tb=12'h845;#1; sino_tb=12'h846;#1; sino_tb=12'h847;#1; sino_tb=12'h848;#1; sino_tb=12'h849;#1; sino_tb=12'h849;#1; sino_tb=12'h84a;#1; 
sino_tb=12'h84b;#1; sino_tb=12'h84c;#1; sino_tb=12'h84d;#1; sino_tb=12'h84e;#1; sino_tb=12'h84f;#1; sino_tb=12'h84f;#1; sino_tb=12'h850;#1; sino_tb=12'h851;#1; 
sino_tb=12'h852;#1; sino_tb=12'h853;#1; sino_tb=12'h854;#1; sino_tb=12'h855;#1; sino_tb=12'h856;#1; sino_tb=12'h856;#1; sino_tb=12'h857;#1; sino_tb=12'h858;#1; 
sino_tb=12'h859;#1; sino_tb=12'h85a;#1; sino_tb=12'h85b;#1; sino_tb=12'h85c;#1; sino_tb=12'h85d;#1; sino_tb=12'h85e;#1; sino_tb=12'h85f;#1; sino_tb=12'h860;#1; 
sino_tb=12'h861;#1; sino_tb=12'h862;#1; sino_tb=12'h862;#1; sino_tb=12'h863;#1; sino_tb=12'h864;#1; sino_tb=12'h865;#1; sino_tb=12'h866;#1; sino_tb=12'h867;#1; 
sino_tb=12'h868;#1; sino_tb=12'h869;#1; sino_tb=12'h86a;#1; sino_tb=12'h86b;#1; sino_tb=12'h86c;#1; sino_tb=12'h86d;#1; sino_tb=12'h86e;#1; sino_tb=12'h86f;#1; 
sino_tb=12'h870;#1; sino_tb=12'h871;#1; sino_tb=12'h872;#1; sino_tb=12'h873;#1; sino_tb=12'h874;#1; sino_tb=12'h876;#1; sino_tb=12'h877;#1; sino_tb=12'h878;#1; 
sino_tb=12'h879;#1; sino_tb=12'h87a;#1; sino_tb=12'h87b;#1; sino_tb=12'h87c;#1; sino_tb=12'h87d;#1; sino_tb=12'h87e;#1; sino_tb=12'h87f;#1; sino_tb=12'h880;#1; 
sino_tb=12'h881;#1; sino_tb=12'h882;#1; sino_tb=12'h883;#1; sino_tb=12'h885;#1; sino_tb=12'h886;#1; sino_tb=12'h887;#1; sino_tb=12'h888;#1; sino_tb=12'h889;#1; 
sino_tb=12'h88a;#1; sino_tb=12'h88b;#1; sino_tb=12'h88c;#1; sino_tb=12'h88e;#1; sino_tb=12'h88f;#1; sino_tb=12'h890;#1; sino_tb=12'h891;#1; sino_tb=12'h892;#1; 
sino_tb=12'h893;#1; sino_tb=12'h895;#1; sino_tb=12'h896;#1; sino_tb=12'h897;#1; sino_tb=12'h898;#1; sino_tb=12'h899;#1; sino_tb=12'h89a;#1; sino_tb=12'h89c;#1; 
sino_tb=12'h89d;#1; sino_tb=12'h89e;#1; sino_tb=12'h89f;#1; sino_tb=12'h8a0;#1; sino_tb=12'h8a2;#1; sino_tb=12'h8a3;#1; sino_tb=12'h8a4;#1; sino_tb=12'h8a5;#1; 
sino_tb=12'h8a7;#1; sino_tb=12'h8a8;#1; sino_tb=12'h8a9;#1; sino_tb=12'h8aa;#1; sino_tb=12'h8ac;#1; sino_tb=12'h8ad;#1; sino_tb=12'h8ae;#1; sino_tb=12'h8af;#1; 
sino_tb=12'h8b1;#1; sino_tb=12'h8b2;#1; sino_tb=12'h8b3;#1; sino_tb=12'h8b4;#1; sino_tb=12'h8b6;#1; sino_tb=12'h8b7;#1; sino_tb=12'h8b8;#1; sino_tb=12'h8ba;#1; 
sino_tb=12'h8bb;#1; sino_tb=12'h8bc;#1; sino_tb=12'h8be;#1; sino_tb=12'h8bf;#1; sino_tb=12'h8c0;#1; sino_tb=12'h8c2;#1; sino_tb=12'h8c3;#1; sino_tb=12'h8c4;#1; 
sino_tb=12'h8c6;#1; sino_tb=12'h8c7;#1; sino_tb=12'h8c8;#1; sino_tb=12'h8ca;#1; sino_tb=12'h8cb;#1; sino_tb=12'h8cc;#1; sino_tb=12'h8ce;#1; sino_tb=12'h8cf;#1; 
sino_tb=12'h8d0;#1; sino_tb=12'h8d2;#1; sino_tb=12'h8d3;#1; sino_tb=12'h8d5;#1; sino_tb=12'h8d6;#1; sino_tb=12'h8d7;#1; sino_tb=12'h8d9;#1; sino_tb=12'h8da;#1; 
sino_tb=12'h8dc;#1; sino_tb=12'h8dd;#1; sino_tb=12'h8de;#1; sino_tb=12'h8e0;#1; sino_tb=12'h8e1;#1; sino_tb=12'h8e3;#1; sino_tb=12'h8e4;#1; sino_tb=12'h8e6;#1; 
sino_tb=12'h8e7;#1; sino_tb=12'h8e8;#1; sino_tb=12'h8ea;#1; sino_tb=12'h8eb;#1; sino_tb=12'h8ed;#1; sino_tb=12'h8ee;#1; sino_tb=12'h8f0;#1; sino_tb=12'h8f1;#1; 
sino_tb=12'h8f3;#1; sino_tb=12'h8f4;#1; sino_tb=12'h8f6;#1; sino_tb=12'h8f7;#1; sino_tb=12'h8f9;#1; sino_tb=12'h8fa;#1; sino_tb=12'h8fc;#1; sino_tb=12'h8fd;#1; 
sino_tb=12'h8ff;#1; sino_tb=12'h900;#1; sino_tb=12'h902;#1; sino_tb=12'h903;#1; sino_tb=12'h905;#1; sino_tb=12'h906;#1; sino_tb=12'h908;#1; sino_tb=12'h909;#1; 
sino_tb=12'h90b;#1; sino_tb=12'h90c;#1; sino_tb=12'h90e;#1; sino_tb=12'h910;#1; sino_tb=12'h911;#1; sino_tb=12'h913;#1; sino_tb=12'h914;#1; sino_tb=12'h916;#1; 
sino_tb=12'h917;#1; sino_tb=12'h919;#1; sino_tb=12'h91b;#1; sino_tb=12'h91c;#1; sino_tb=12'h91e;#1; sino_tb=12'h91f;#1; sino_tb=12'h921;#1; sino_tb=12'h923;#1; 
sino_tb=12'h924;#1; sino_tb=12'h926;#1; sino_tb=12'h927;#1; sino_tb=12'h929;#1; sino_tb=12'h92b;#1; sino_tb=12'h92c;#1; sino_tb=12'h92e;#1; sino_tb=12'h930;#1; 
sino_tb=12'h931;#1; sino_tb=12'h933;#1; sino_tb=12'h935;#1; sino_tb=12'h936;#1; sino_tb=12'h938;#1; sino_tb=12'h93a;#1; sino_tb=12'h93b;#1; sino_tb=12'h93d;#1; 
sino_tb=12'h93f;#1; sino_tb=12'h940;#1; sino_tb=12'h942;#1; sino_tb=12'h944;#1; sino_tb=12'h945;#1; sino_tb=12'h947;#1; sino_tb=12'h949;#1; sino_tb=12'h94a;#1; 
sino_tb=12'h94c;#1; sino_tb=12'h94e;#1; sino_tb=12'h950;#1; sino_tb=12'h951;#1; sino_tb=12'h953;#1; sino_tb=12'h955;#1; sino_tb=12'h957;#1; sino_tb=12'h958;#1; 
sino_tb=12'h95a;#1; sino_tb=12'h95c;#1; sino_tb=12'h95d;#1; sino_tb=12'h95f;#1; sino_tb=12'h961;#1; sino_tb=12'h963;#1; sino_tb=12'h965;#1; sino_tb=12'h966;#1; 
sino_tb=12'h968;#1; sino_tb=12'h96a;#1; sino_tb=12'h96c;#1; sino_tb=12'h96d;#1; sino_tb=12'h96f;#1; sino_tb=12'h971;#1; sino_tb=12'h973;#1; sino_tb=12'h975;#1; 
sino_tb=12'h976;#1; sino_tb=12'h978;#1; sino_tb=12'h97a;#1; sino_tb=12'h97c;#1; sino_tb=12'h97e;#1; sino_tb=12'h97f;#1; sino_tb=12'h981;#1; sino_tb=12'h983;#1; 
sino_tb=12'h985;#1; sino_tb=12'h987;#1; sino_tb=12'h989;#1; sino_tb=12'h98b;#1; sino_tb=12'h98c;#1; sino_tb=12'h98e;#1; sino_tb=12'h990;#1; sino_tb=12'h992;#1; 
sino_tb=12'h994;#1; sino_tb=12'h996;#1; sino_tb=12'h998;#1; sino_tb=12'h999;#1; sino_tb=12'h99b;#1; sino_tb=12'h99d;#1; sino_tb=12'h99f;#1; sino_tb=12'h9a1;#1; 
sino_tb=12'h9a3;#1; sino_tb=12'h9a5;#1; sino_tb=12'h9a7;#1; sino_tb=12'h9a9;#1; sino_tb=12'h9ab;#1; sino_tb=12'h9ac;#1; sino_tb=12'h9ae;#1; sino_tb=12'h9b0;#1; 
sino_tb=12'h9b2;#1; sino_tb=12'h9b4;#1; sino_tb=12'h9b6;#1; sino_tb=12'h9b8;#1; sino_tb=12'h9ba;#1; sino_tb=12'h9bc;#1; sino_tb=12'h9be;#1; sino_tb=12'h9c0;#1; 
sino_tb=12'h9c2;#1; sino_tb=12'h9c4;#1; sino_tb=12'h9c6;#1; sino_tb=12'h9c8;#1; sino_tb=12'h9ca;#1; sino_tb=12'h9cc;#1; sino_tb=12'h9ce;#1; sino_tb=12'h9d0;#1; 
sino_tb=12'h9d2;#1; sino_tb=12'h9d4;#1; sino_tb=12'h9d6;#1; sino_tb=12'h9d8;#1; sino_tb=12'h9da;#1; sino_tb=12'h9dc;#1; sino_tb=12'h9de;#1; sino_tb=12'h9e0;#1; 
sino_tb=12'h9e2;#1; sino_tb=12'h9e4;#1; sino_tb=12'h9e6;#1; sino_tb=12'h9e8;#1; sino_tb=12'h9ea;#1; sino_tb=12'h9ec;#1; sino_tb=12'h9ee;#1; sino_tb=12'h9f0;#1; 
sino_tb=12'h9f2;#1; sino_tb=12'h9f4;#1; sino_tb=12'h9f6;#1; sino_tb=12'h9f8;#1; sino_tb=12'h9fa;#1; sino_tb=12'h9fc;#1; sino_tb=12'h9fe;#1; sino_tb=12'ha00;#1; 
sino_tb=12'ha03;#1; sino_tb=12'ha05;#1; sino_tb=12'ha07;#1; sino_tb=12'ha09;#1; sino_tb=12'ha0b;#1; sino_tb=12'ha0d;#1; sino_tb=12'ha0f;#1; sino_tb=12'ha11;#1; 
sino_tb=12'ha13;#1; sino_tb=12'ha15;#1; sino_tb=12'ha17;#1; sino_tb=12'ha1a;#1; sino_tb=12'ha1c;#1; sino_tb=12'ha1e;#1; sino_tb=12'ha20;#1; sino_tb=12'ha22;#1; 
sino_tb=12'ha24;#1; sino_tb=12'ha26;#1; sino_tb=12'ha29;#1; sino_tb=12'ha2b;#1; sino_tb=12'ha2d;#1; sino_tb=12'ha2f;#1; sino_tb=12'ha31;#1; sino_tb=12'ha33;#1; 
sino_tb=12'ha35;#1; sino_tb=12'ha38;#1; sino_tb=12'ha3a;#1; sino_tb=12'ha3c;#1; sino_tb=12'ha3e;#1; sino_tb=12'ha40;#1; sino_tb=12'ha43;#1; sino_tb=12'ha45;#1; 
sino_tb=12'ha47;#1; sino_tb=12'ha49;#1; sino_tb=12'ha4b;#1; sino_tb=12'ha4d;#1; sino_tb=12'ha50;#1; sino_tb=12'ha52;#1; sino_tb=12'ha54;#1; sino_tb=12'ha56;#1; 
sino_tb=12'ha59;#1; sino_tb=12'ha5b;#1; sino_tb=12'ha5d;#1; sino_tb=12'ha5f;#1; sino_tb=12'ha61;#1; sino_tb=12'ha64;#1; sino_tb=12'ha66;#1; sino_tb=12'ha68;#1; 
sino_tb=12'ha6a;#1; sino_tb=12'ha6d;#1; sino_tb=12'ha6f;#1; sino_tb=12'ha71;#1; sino_tb=12'ha73;#1; sino_tb=12'ha76;#1; sino_tb=12'ha78;#1; sino_tb=12'ha7a;#1; 
sino_tb=12'ha7d;#1; sino_tb=12'ha7f;#1; sino_tb=12'ha81;#1; sino_tb=12'ha83;#1; sino_tb=12'ha86;#1; sino_tb=12'ha88;#1; sino_tb=12'ha8a;#1; sino_tb=12'ha8d;#1; 
sino_tb=12'ha8f;#1; sino_tb=12'ha91;#1; sino_tb=12'ha93;#1; sino_tb=12'ha96;#1; sino_tb=12'ha98;#1; sino_tb=12'ha9a;#1; sino_tb=12'ha9d;#1; sino_tb=12'ha9f;#1; 
sino_tb=12'haa1;#1; sino_tb=12'haa4;#1; sino_tb=12'haa6;#1; sino_tb=12'haa8;#1; sino_tb=12'haab;#1; sino_tb=12'haad;#1; sino_tb=12'haaf;#1; sino_tb=12'hab2;#1; 
sino_tb=12'hab4;#1; sino_tb=12'hab6;#1; sino_tb=12'hab9;#1; sino_tb=12'habb;#1; sino_tb=12'habd;#1; sino_tb=12'hac0;#1; sino_tb=12'hac2;#1; sino_tb=12'hac5;#1; 
sino_tb=12'hac7;#1; sino_tb=12'hac9;#1; sino_tb=12'hacc;#1; sino_tb=12'hace;#1; sino_tb=12'had0;#1; sino_tb=12'had3;#1; sino_tb=12'had5;#1; sino_tb=12'had8;#1; 
sino_tb=12'hada;#1; sino_tb=12'hadc;#1; sino_tb=12'hadf;#1; sino_tb=12'hae1;#1; sino_tb=12'hae4;#1; sino_tb=12'hae6;#1; sino_tb=12'hae9;#1; sino_tb=12'haeb;#1; 
sino_tb=12'haed;#1; sino_tb=12'haf0;#1; sino_tb=12'haf2;#1; sino_tb=12'haf5;#1; sino_tb=12'haf7;#1; sino_tb=12'hafa;#1; sino_tb=12'hafc;#1; sino_tb=12'hafe;#1; 
sino_tb=12'hb01;#1; sino_tb=12'hb03;#1; sino_tb=12'hb06;#1; sino_tb=12'hb08;#1; sino_tb=12'hb0b;#1; sino_tb=12'hb0d;#1; sino_tb=12'hb10;#1; sino_tb=12'hb12;#1; 
sino_tb=12'hb15;#1; sino_tb=12'hb17;#1; sino_tb=12'hb1a;#1; sino_tb=12'hb1c;#1; sino_tb=12'hb1f;#1; sino_tb=12'hb21;#1; sino_tb=12'hb24;#1; sino_tb=12'hb26;#1; 
sino_tb=12'hb29;#1; sino_tb=12'hb2b;#1; sino_tb=12'hb2e;#1; sino_tb=12'hb30;#1; sino_tb=12'hb33;#1; sino_tb=12'hb35;#1; sino_tb=12'hb38;#1; sino_tb=12'hb3a;#1; 
sino_tb=12'hb3d;#1; sino_tb=12'hb3f;#1; sino_tb=12'hb42;#1; sino_tb=12'hb44;#1; sino_tb=12'hb47;#1; sino_tb=12'hb49;#1; sino_tb=12'hb4c;#1; sino_tb=12'hb4e;#1; 
sino_tb=12'hb51;#1; sino_tb=12'hb53;#1; sino_tb=12'hb56;#1; sino_tb=12'hb59;#1; sino_tb=12'hb5b;#1; sino_tb=12'hb5e;#1; sino_tb=12'hb60;#1; sino_tb=12'hb63;#1; 
sino_tb=12'hb65;#1; sino_tb=12'hb68;#1; sino_tb=12'hb6a;#1; sino_tb=12'hb6d;#1; sino_tb=12'hb70;#1; sino_tb=12'hb72;#1; sino_tb=12'hb75;#1; sino_tb=12'hb77;#1; 
sino_tb=12'hb7a;#1; sino_tb=12'hb7d;#1; sino_tb=12'hb7f;#1; sino_tb=12'hb82;#1; sino_tb=12'hb84;#1; sino_tb=12'hb87;#1; sino_tb=12'hb8a;#1; sino_tb=12'hb8c;#1; 
sino_tb=12'hb8f;#1; sino_tb=12'hb91;#1; sino_tb=12'hb94;#1; sino_tb=12'hb97;#1; sino_tb=12'hb99;#1; sino_tb=12'hb9c;#1; sino_tb=12'hb9e;#1; sino_tb=12'hba1;#1; 
sino_tb=12'hba4;#1; sino_tb=12'hba6;#1; sino_tb=12'hba9;#1; sino_tb=12'hbac;#1; sino_tb=12'hbae;#1; sino_tb=12'hbb1;#1; sino_tb=12'hbb4;#1; sino_tb=12'hbb6;#1; 
sino_tb=12'hbb9;#1; sino_tb=12'hbbc;#1; sino_tb=12'hbbe;#1; sino_tb=12'hbc1;#1; sino_tb=12'hbc3;#1; sino_tb=12'hbc6;#1; sino_tb=12'hbc9;#1; sino_tb=12'hbcb;#1; 
sino_tb=12'hbce;#1; sino_tb=12'hbd1;#1; sino_tb=12'hbd4;#1; sino_tb=12'hbd6;#1; sino_tb=12'hbd9;#1; sino_tb=12'hbdc;#1; sino_tb=12'hbde;#1; sino_tb=12'hbe1;#1; 
sino_tb=12'hbe4;#1; sino_tb=12'hbe6;#1; sino_tb=12'hbe9;#1; sino_tb=12'hbec;#1; sino_tb=12'hbee;#1; sino_tb=12'hbf1;#1; sino_tb=12'hbf4;#1; sino_tb=12'hbf7;#1; 
sino_tb=12'hbf9;#1; sino_tb=12'hbfc;#1; sino_tb=12'hbff;#1; sino_tb=12'hc01;#1; sino_tb=12'hc04;#1; sino_tb=12'hc07;#1; sino_tb=12'hc0a;#1; sino_tb=12'hc0c;#1; 
sino_tb=12'hc0f;#1; sino_tb=12'hc12;#1; sino_tb=12'hc15;#1; sino_tb=12'hc17;#1; sino_tb=12'hc1a;#1; sino_tb=12'hc1d;#1; sino_tb=12'hc1f;#1; sino_tb=12'hc22;#1; 
sino_tb=12'hc25;#1; sino_tb=12'hc28;#1; sino_tb=12'hc2a;#1; sino_tb=12'hc2d;#1; sino_tb=12'hc30;#1; sino_tb=12'hc33;#1; sino_tb=12'hc36;#1; sino_tb=12'hc38;#1; 
sino_tb=12'hc3b;#1; sino_tb=12'hc3e;#1; sino_tb=12'hc41;#1; sino_tb=12'hc43;#1; sino_tb=12'hc46;#1; sino_tb=12'hc49;#1; sino_tb=12'hc4c;#1; sino_tb=12'hc4e;#1; 
sino_tb=12'hc51;#1; sino_tb=12'hc54;#1; sino_tb=12'hc57;#1; sino_tb=12'hc5a;#1; sino_tb=12'hc5c;#1; sino_tb=12'hc5f;#1; sino_tb=12'hc62;#1; sino_tb=12'hc65;#1; 
sino_tb=12'hc68;#1; sino_tb=12'hc6a;#1; sino_tb=12'hc6d;#1; sino_tb=12'hc70;#1; sino_tb=12'hc73;#1; sino_tb=12'hc76;#1; sino_tb=12'hc79;#1; sino_tb=12'hc7b;#1; 
sino_tb=12'hc7e;#1; sino_tb=12'hc81;#1; sino_tb=12'hc84;#1; sino_tb=12'hc87;#1; sino_tb=12'hc89;#1; sino_tb=12'hc8c;#1; sino_tb=12'hc8f;#1; sino_tb=12'hc92;#1; 
sino_tb=12'hc95;#1; sino_tb=12'hc98;#1; sino_tb=12'hc9a;#1; sino_tb=12'hc9d;#1; sino_tb=12'hca0;#1; sino_tb=12'hca3;#1; sino_tb=12'hca6;#1; sino_tb=12'hca9;#1; 
sino_tb=12'hcac;#1; sino_tb=12'hcae;#1; sino_tb=12'hcb1;#1; sino_tb=12'hcb4;#1; sino_tb=12'hcb7;#1; sino_tb=12'hcba;#1; sino_tb=12'hcbd;#1; sino_tb=12'hcc0;#1; 
sino_tb=12'hcc2;#1; sino_tb=12'hcc5;#1; sino_tb=12'hcc8;#1; sino_tb=12'hccb;#1; sino_tb=12'hcce;#1; sino_tb=12'hcd1;#1; sino_tb=12'hcd4;#1; sino_tb=12'hcd7;#1; 
sino_tb=12'hcd9;#1; sino_tb=12'hcdc;#1; sino_tb=12'hcdf;#1; sino_tb=12'hce2;#1; sino_tb=12'hce5;#1; sino_tb=12'hce8;#1; sino_tb=12'hceb;#1; sino_tb=12'hcee;#1; 
sino_tb=12'hcf1;#1; sino_tb=12'hcf4;#1; sino_tb=12'hcf6;#1; sino_tb=12'hcf9;#1; sino_tb=12'hcfc;#1; sino_tb=12'hcff;#1; sino_tb=12'hd02;#1; sino_tb=12'hd05;#1; 
sino_tb=12'hd08;#1; sino_tb=12'hd0b;#1; sino_tb=12'hd0e;#1; sino_tb=12'hd11;#1; sino_tb=12'hd14;#1; sino_tb=12'hd17;#1; sino_tb=12'hd19;#1; sino_tb=12'hd1c;#1; 
sino_tb=12'hd1f;#1; sino_tb=12'hd22;#1; sino_tb=12'hd25;#1; sino_tb=12'hd28;#1; sino_tb=12'hd2b;#1; sino_tb=12'hd2e;#1; sino_tb=12'hd31;#1; sino_tb=12'hd34;#1; 
sino_tb=12'hd37;#1; sino_tb=12'hd3a;#1; sino_tb=12'hd3d;#1; sino_tb=12'hd40;#1; sino_tb=12'hd43;#1; sino_tb=12'hd46;#1; sino_tb=12'hd48;#1; sino_tb=12'hd4b;#1; 
sino_tb=12'hd4e;#1; sino_tb=12'hd51;#1; sino_tb=12'hd54;#1; sino_tb=12'hd57;#1; sino_tb=12'hd5a;#1; sino_tb=12'hd5d;#1; sino_tb=12'hd60;#1; sino_tb=12'hd63;#1; 
sino_tb=12'hd66;#1; sino_tb=12'hd69;#1; sino_tb=12'hd6c;#1; sino_tb=12'hd6f;#1; sino_tb=12'hd72;#1; sino_tb=12'hd75;#1; sino_tb=12'hd78;#1; sino_tb=12'hd7b;#1; 
sino_tb=12'hd7e;#1; sino_tb=12'hd81;#1; sino_tb=12'hd84;#1; sino_tb=12'hd87;#1; sino_tb=12'hd8a;#1; sino_tb=12'hd8d;#1; sino_tb=12'hd90;#1; sino_tb=12'hd93;#1; 
sino_tb=12'hd96;#1; sino_tb=12'hd99;#1; sino_tb=12'hd9c;#1; sino_tb=12'hd9f;#1; sino_tb=12'hda2;#1; sino_tb=12'hda5;#1; sino_tb=12'hda8;#1; sino_tb=12'hdab;#1; 
sino_tb=12'hdae;#1; sino_tb=12'hdb1;#1; sino_tb=12'hdb4;#1; sino_tb=12'hdb7;#1; sino_tb=12'hdba;#1; sino_tb=12'hdbd;#1; sino_tb=12'hdc0;#1; sino_tb=12'hdc3;#1; 
sino_tb=12'hdc6;#1; sino_tb=12'hdc9;#1; sino_tb=12'hdcc;#1; sino_tb=12'hdcf;#1; sino_tb=12'hdd2;#1; sino_tb=12'hdd5;#1; sino_tb=12'hdd8;#1; sino_tb=12'hddb;#1; 
sino_tb=12'hdde;#1; sino_tb=12'hde1;#1; sino_tb=12'hde4;#1; sino_tb=12'hde7;#1; sino_tb=12'hdea;#1; sino_tb=12'hded;#1; sino_tb=12'hdf0;#1; sino_tb=12'hdf3;#1; 
sino_tb=12'hdf6;#1; sino_tb=12'hdf9;#1; sino_tb=12'hdfc;#1; sino_tb=12'hdff;#1; sino_tb=12'he02;#1; sino_tb=12'he05;#1; sino_tb=12'he09;#1; sino_tb=12'he0c;#1; 
sino_tb=12'he0f;#1; sino_tb=12'he12;#1; sino_tb=12'he15;#1; sino_tb=12'he18;#1; sino_tb=12'he1b;#1; sino_tb=12'he1e;#1; sino_tb=12'he21;#1; sino_tb=12'he24;#1; 
sino_tb=12'he27;#1; sino_tb=12'he2a;#1; sino_tb=12'he2d;#1; sino_tb=12'he30;#1; sino_tb=12'he33;#1; sino_tb=12'he36;#1; sino_tb=12'he39;#1; sino_tb=12'he3c;#1; 
sino_tb=12'he3f;#1; sino_tb=12'he43;#1; sino_tb=12'he46;#1; sino_tb=12'he49;#1; sino_tb=12'he4c;#1; sino_tb=12'he4f;#1; sino_tb=12'he52;#1; sino_tb=12'he55;#1; 
sino_tb=12'he58;#1; sino_tb=12'he5b;#1; sino_tb=12'he5e;#1; sino_tb=12'he61;#1; sino_tb=12'he64;#1; sino_tb=12'he67;#1; sino_tb=12'he6a;#1; sino_tb=12'he6e;#1; 
sino_tb=12'he71;#1; sino_tb=12'he74;#1; sino_tb=12'he77;#1; sino_tb=12'he7a;#1; sino_tb=12'he7d;#1; sino_tb=12'he80;#1; sino_tb=12'he83;#1; sino_tb=12'he86;#1; 
sino_tb=12'he89;#1; sino_tb=12'he8c;#1; sino_tb=12'he8f;#1; sino_tb=12'he93;#1; sino_tb=12'he96;#1; sino_tb=12'he99;#1; sino_tb=12'he9c;#1; sino_tb=12'he9f;#1; 
sino_tb=12'hea2;#1; sino_tb=12'hea5;#1; sino_tb=12'hea8;#1; sino_tb=12'heab;#1; sino_tb=12'heae;#1; sino_tb=12'heb2;#1; sino_tb=12'heb5;#1; sino_tb=12'heb8;#1; 
sino_tb=12'hebb;#1; sino_tb=12'hebe;#1; sino_tb=12'hec1;#1; sino_tb=12'hec4;#1; sino_tb=12'hec7;#1; sino_tb=12'heca;#1; sino_tb=12'hecd;#1; sino_tb=12'hed1;#1; 
sino_tb=12'hed4;#1; sino_tb=12'hed7;#1; sino_tb=12'heda;#1; sino_tb=12'hedd;#1; sino_tb=12'hee0;#1; sino_tb=12'hee3;#1; sino_tb=12'hee6;#1; sino_tb=12'hee9;#1; 
sino_tb=12'heed;#1; sino_tb=12'hef0;#1; sino_tb=12'hef3;#1; sino_tb=12'hef6;#1; sino_tb=12'hef9;#1; sino_tb=12'hefc;#1; sino_tb=12'heff;#1; sino_tb=12'hf02;#1; 
sino_tb=12'hf05;#1; sino_tb=12'hf09;#1; sino_tb=12'hf0c;#1; sino_tb=12'hf0f;#1; sino_tb=12'hf12;#1; sino_tb=12'hf15;#1; sino_tb=12'hf18;#1; sino_tb=12'hf1b;#1; 
sino_tb=12'hf1e;#1; sino_tb=12'hf21;#1; sino_tb=12'hf25;#1; sino_tb=12'hf28;#1; sino_tb=12'hf2b;#1; sino_tb=12'hf2e;#1; sino_tb=12'hf31;#1; sino_tb=12'hf34;#1; 
sino_tb=12'hf37;#1; sino_tb=12'hf3a;#1; sino_tb=12'hf3e;#1; sino_tb=12'hf41;#1; sino_tb=12'hf44;#1; sino_tb=12'hf47;#1; sino_tb=12'hf4a;#1; sino_tb=12'hf4d;#1; 
sino_tb=12'hf50;#1; sino_tb=12'hf54;#1; sino_tb=12'hf57;#1; sino_tb=12'hf5a;#1; sino_tb=12'hf5d;#1; sino_tb=12'hf60;#1; sino_tb=12'hf63;#1; sino_tb=12'hf66;#1; 
sino_tb=12'hf69;#1; sino_tb=12'hf6d;#1; sino_tb=12'hf70;#1; sino_tb=12'hf73;#1; sino_tb=12'hf76;#1; sino_tb=12'hf79;#1; sino_tb=12'hf7c;#1; sino_tb=12'hf7f;#1; 
sino_tb=12'hf82;#1; sino_tb=12'hf86;#1; sino_tb=12'hf89;#1; sino_tb=12'hf8c;#1; sino_tb=12'hf8f;#1; sino_tb=12'hf92;#1; sino_tb=12'hf95;#1; sino_tb=12'hf98;#1; 
sino_tb=12'hf9c;#1; sino_tb=12'hf9f;#1; sino_tb=12'hfa2;#1; sino_tb=12'hfa5;#1; sino_tb=12'hfa8;#1; sino_tb=12'hfab;#1; sino_tb=12'hfae;#1; sino_tb=12'hfb2;#1; 
sino_tb=12'hfb5;#1; sino_tb=12'hfb8;#1; sino_tb=12'hfbb;#1; sino_tb=12'hfbe;#1; sino_tb=12'hfc1;#1; sino_tb=12'hfc4;#1; sino_tb=12'hfc7;#1; sino_tb=12'hfcb;#1; 
sino_tb=12'hfce;#1; sino_tb=12'hfd1;#1; sino_tb=12'hfd4;#1; sino_tb=12'hfd7;#1; sino_tb=12'hfda;#1; sino_tb=12'hfdd;#1; sino_tb=12'hfe1;#1; sino_tb=12'hfe4;#1; 
sino_tb=12'hfe7;#1; sino_tb=12'hfea;#1; sino_tb=12'hfed;#1; sino_tb=12'hff0;#1; sino_tb=12'hff3;#1; sino_tb=12'hff7;#1; sino_tb=12'hffa;#1; sino_tb=12'hffd;


end


endmodule