module key_search();


endmodule