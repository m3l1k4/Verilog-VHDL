module test();


always@(posedge clk) begin


end 

endmodule