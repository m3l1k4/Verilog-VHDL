module loop_3(
input logic clk,
input logic reset,
input logic start_flag,
input logic [7:0] data_in,
output logic [7:0] data_out,



); 



endmodule 